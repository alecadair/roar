MACRO NMOS_S_65192303_X16_Y6
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_65192303_X16_Y6 0 0 ;
  SIZE 15480 BY 36960 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 7170 260 7450 29980 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 7600 4460 7880 34180 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 8030 680 8310 36280 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 36625 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 33265 ;
    LAYER M1 ;
      RECT 2025 33515 2275 34525 ;
    LAYER M1 ;
      RECT 2025 35615 2275 36625 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 15625 ;
    LAYER M1 ;
      RECT 2885 15875 3135 16885 ;
    LAYER M1 ;
      RECT 2885 17975 3135 21505 ;
    LAYER M1 ;
      RECT 2885 21755 3135 22765 ;
    LAYER M1 ;
      RECT 2885 23855 3135 27385 ;
    LAYER M1 ;
      RECT 2885 27635 3135 28645 ;
    LAYER M1 ;
      RECT 2885 29735 3135 33265 ;
    LAYER M1 ;
      RECT 2885 33515 3135 34525 ;
    LAYER M1 ;
      RECT 2885 35615 3135 36625 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 23855 3565 27385 ;
    LAYER M1 ;
      RECT 3315 29735 3565 33265 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 15625 ;
    LAYER M1 ;
      RECT 3745 15875 3995 16885 ;
    LAYER M1 ;
      RECT 3745 17975 3995 21505 ;
    LAYER M1 ;
      RECT 3745 21755 3995 22765 ;
    LAYER M1 ;
      RECT 3745 23855 3995 27385 ;
    LAYER M1 ;
      RECT 3745 27635 3995 28645 ;
    LAYER M1 ;
      RECT 3745 29735 3995 33265 ;
    LAYER M1 ;
      RECT 3745 33515 3995 34525 ;
    LAYER M1 ;
      RECT 3745 35615 3995 36625 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4175 17975 4425 21505 ;
    LAYER M1 ;
      RECT 4175 23855 4425 27385 ;
    LAYER M1 ;
      RECT 4175 29735 4425 33265 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 15625 ;
    LAYER M1 ;
      RECT 4605 15875 4855 16885 ;
    LAYER M1 ;
      RECT 4605 17975 4855 21505 ;
    LAYER M1 ;
      RECT 4605 21755 4855 22765 ;
    LAYER M1 ;
      RECT 4605 23855 4855 27385 ;
    LAYER M1 ;
      RECT 4605 27635 4855 28645 ;
    LAYER M1 ;
      RECT 4605 29735 4855 33265 ;
    LAYER M1 ;
      RECT 4605 33515 4855 34525 ;
    LAYER M1 ;
      RECT 4605 35615 4855 36625 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5035 12095 5285 15625 ;
    LAYER M1 ;
      RECT 5035 17975 5285 21505 ;
    LAYER M1 ;
      RECT 5035 23855 5285 27385 ;
    LAYER M1 ;
      RECT 5035 29735 5285 33265 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 15625 ;
    LAYER M1 ;
      RECT 5465 15875 5715 16885 ;
    LAYER M1 ;
      RECT 5465 17975 5715 21505 ;
    LAYER M1 ;
      RECT 5465 21755 5715 22765 ;
    LAYER M1 ;
      RECT 5465 23855 5715 27385 ;
    LAYER M1 ;
      RECT 5465 27635 5715 28645 ;
    LAYER M1 ;
      RECT 5465 29735 5715 33265 ;
    LAYER M1 ;
      RECT 5465 33515 5715 34525 ;
    LAYER M1 ;
      RECT 5465 35615 5715 36625 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 5895 12095 6145 15625 ;
    LAYER M1 ;
      RECT 5895 17975 6145 21505 ;
    LAYER M1 ;
      RECT 5895 23855 6145 27385 ;
    LAYER M1 ;
      RECT 5895 29735 6145 33265 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 9745 ;
    LAYER M1 ;
      RECT 6325 9995 6575 11005 ;
    LAYER M1 ;
      RECT 6325 12095 6575 15625 ;
    LAYER M1 ;
      RECT 6325 15875 6575 16885 ;
    LAYER M1 ;
      RECT 6325 17975 6575 21505 ;
    LAYER M1 ;
      RECT 6325 21755 6575 22765 ;
    LAYER M1 ;
      RECT 6325 23855 6575 27385 ;
    LAYER M1 ;
      RECT 6325 27635 6575 28645 ;
    LAYER M1 ;
      RECT 6325 29735 6575 33265 ;
    LAYER M1 ;
      RECT 6325 33515 6575 34525 ;
    LAYER M1 ;
      RECT 6325 35615 6575 36625 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 6215 7005 9745 ;
    LAYER M1 ;
      RECT 6755 12095 7005 15625 ;
    LAYER M1 ;
      RECT 6755 17975 7005 21505 ;
    LAYER M1 ;
      RECT 6755 23855 7005 27385 ;
    LAYER M1 ;
      RECT 6755 29735 7005 33265 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 9745 ;
    LAYER M1 ;
      RECT 7185 9995 7435 11005 ;
    LAYER M1 ;
      RECT 7185 12095 7435 15625 ;
    LAYER M1 ;
      RECT 7185 15875 7435 16885 ;
    LAYER M1 ;
      RECT 7185 17975 7435 21505 ;
    LAYER M1 ;
      RECT 7185 21755 7435 22765 ;
    LAYER M1 ;
      RECT 7185 23855 7435 27385 ;
    LAYER M1 ;
      RECT 7185 27635 7435 28645 ;
    LAYER M1 ;
      RECT 7185 29735 7435 33265 ;
    LAYER M1 ;
      RECT 7185 33515 7435 34525 ;
    LAYER M1 ;
      RECT 7185 35615 7435 36625 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 7615 6215 7865 9745 ;
    LAYER M1 ;
      RECT 7615 12095 7865 15625 ;
    LAYER M1 ;
      RECT 7615 17975 7865 21505 ;
    LAYER M1 ;
      RECT 7615 23855 7865 27385 ;
    LAYER M1 ;
      RECT 7615 29735 7865 33265 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 9745 ;
    LAYER M1 ;
      RECT 8045 9995 8295 11005 ;
    LAYER M1 ;
      RECT 8045 12095 8295 15625 ;
    LAYER M1 ;
      RECT 8045 15875 8295 16885 ;
    LAYER M1 ;
      RECT 8045 17975 8295 21505 ;
    LAYER M1 ;
      RECT 8045 21755 8295 22765 ;
    LAYER M1 ;
      RECT 8045 23855 8295 27385 ;
    LAYER M1 ;
      RECT 8045 27635 8295 28645 ;
    LAYER M1 ;
      RECT 8045 29735 8295 33265 ;
    LAYER M1 ;
      RECT 8045 33515 8295 34525 ;
    LAYER M1 ;
      RECT 8045 35615 8295 36625 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8475 6215 8725 9745 ;
    LAYER M1 ;
      RECT 8475 12095 8725 15625 ;
    LAYER M1 ;
      RECT 8475 17975 8725 21505 ;
    LAYER M1 ;
      RECT 8475 23855 8725 27385 ;
    LAYER M1 ;
      RECT 8475 29735 8725 33265 ;
    LAYER M1 ;
      RECT 8905 335 9155 3865 ;
    LAYER M1 ;
      RECT 8905 4115 9155 5125 ;
    LAYER M1 ;
      RECT 8905 6215 9155 9745 ;
    LAYER M1 ;
      RECT 8905 9995 9155 11005 ;
    LAYER M1 ;
      RECT 8905 12095 9155 15625 ;
    LAYER M1 ;
      RECT 8905 15875 9155 16885 ;
    LAYER M1 ;
      RECT 8905 17975 9155 21505 ;
    LAYER M1 ;
      RECT 8905 21755 9155 22765 ;
    LAYER M1 ;
      RECT 8905 23855 9155 27385 ;
    LAYER M1 ;
      RECT 8905 27635 9155 28645 ;
    LAYER M1 ;
      RECT 8905 29735 9155 33265 ;
    LAYER M1 ;
      RECT 8905 33515 9155 34525 ;
    LAYER M1 ;
      RECT 8905 35615 9155 36625 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 9335 6215 9585 9745 ;
    LAYER M1 ;
      RECT 9335 12095 9585 15625 ;
    LAYER M1 ;
      RECT 9335 17975 9585 21505 ;
    LAYER M1 ;
      RECT 9335 23855 9585 27385 ;
    LAYER M1 ;
      RECT 9335 29735 9585 33265 ;
    LAYER M1 ;
      RECT 9765 335 10015 3865 ;
    LAYER M1 ;
      RECT 9765 4115 10015 5125 ;
    LAYER M1 ;
      RECT 9765 6215 10015 9745 ;
    LAYER M1 ;
      RECT 9765 9995 10015 11005 ;
    LAYER M1 ;
      RECT 9765 12095 10015 15625 ;
    LAYER M1 ;
      RECT 9765 15875 10015 16885 ;
    LAYER M1 ;
      RECT 9765 17975 10015 21505 ;
    LAYER M1 ;
      RECT 9765 21755 10015 22765 ;
    LAYER M1 ;
      RECT 9765 23855 10015 27385 ;
    LAYER M1 ;
      RECT 9765 27635 10015 28645 ;
    LAYER M1 ;
      RECT 9765 29735 10015 33265 ;
    LAYER M1 ;
      RECT 9765 33515 10015 34525 ;
    LAYER M1 ;
      RECT 9765 35615 10015 36625 ;
    LAYER M1 ;
      RECT 10195 335 10445 3865 ;
    LAYER M1 ;
      RECT 10195 6215 10445 9745 ;
    LAYER M1 ;
      RECT 10195 12095 10445 15625 ;
    LAYER M1 ;
      RECT 10195 17975 10445 21505 ;
    LAYER M1 ;
      RECT 10195 23855 10445 27385 ;
    LAYER M1 ;
      RECT 10195 29735 10445 33265 ;
    LAYER M1 ;
      RECT 10625 335 10875 3865 ;
    LAYER M1 ;
      RECT 10625 4115 10875 5125 ;
    LAYER M1 ;
      RECT 10625 6215 10875 9745 ;
    LAYER M1 ;
      RECT 10625 9995 10875 11005 ;
    LAYER M1 ;
      RECT 10625 12095 10875 15625 ;
    LAYER M1 ;
      RECT 10625 15875 10875 16885 ;
    LAYER M1 ;
      RECT 10625 17975 10875 21505 ;
    LAYER M1 ;
      RECT 10625 21755 10875 22765 ;
    LAYER M1 ;
      RECT 10625 23855 10875 27385 ;
    LAYER M1 ;
      RECT 10625 27635 10875 28645 ;
    LAYER M1 ;
      RECT 10625 29735 10875 33265 ;
    LAYER M1 ;
      RECT 10625 33515 10875 34525 ;
    LAYER M1 ;
      RECT 10625 35615 10875 36625 ;
    LAYER M1 ;
      RECT 11055 335 11305 3865 ;
    LAYER M1 ;
      RECT 11055 6215 11305 9745 ;
    LAYER M1 ;
      RECT 11055 12095 11305 15625 ;
    LAYER M1 ;
      RECT 11055 17975 11305 21505 ;
    LAYER M1 ;
      RECT 11055 23855 11305 27385 ;
    LAYER M1 ;
      RECT 11055 29735 11305 33265 ;
    LAYER M1 ;
      RECT 11485 335 11735 3865 ;
    LAYER M1 ;
      RECT 11485 4115 11735 5125 ;
    LAYER M1 ;
      RECT 11485 6215 11735 9745 ;
    LAYER M1 ;
      RECT 11485 9995 11735 11005 ;
    LAYER M1 ;
      RECT 11485 12095 11735 15625 ;
    LAYER M1 ;
      RECT 11485 15875 11735 16885 ;
    LAYER M1 ;
      RECT 11485 17975 11735 21505 ;
    LAYER M1 ;
      RECT 11485 21755 11735 22765 ;
    LAYER M1 ;
      RECT 11485 23855 11735 27385 ;
    LAYER M1 ;
      RECT 11485 27635 11735 28645 ;
    LAYER M1 ;
      RECT 11485 29735 11735 33265 ;
    LAYER M1 ;
      RECT 11485 33515 11735 34525 ;
    LAYER M1 ;
      RECT 11485 35615 11735 36625 ;
    LAYER M1 ;
      RECT 11915 335 12165 3865 ;
    LAYER M1 ;
      RECT 11915 6215 12165 9745 ;
    LAYER M1 ;
      RECT 11915 12095 12165 15625 ;
    LAYER M1 ;
      RECT 11915 17975 12165 21505 ;
    LAYER M1 ;
      RECT 11915 23855 12165 27385 ;
    LAYER M1 ;
      RECT 11915 29735 12165 33265 ;
    LAYER M1 ;
      RECT 12345 335 12595 3865 ;
    LAYER M1 ;
      RECT 12345 4115 12595 5125 ;
    LAYER M1 ;
      RECT 12345 6215 12595 9745 ;
    LAYER M1 ;
      RECT 12345 9995 12595 11005 ;
    LAYER M1 ;
      RECT 12345 12095 12595 15625 ;
    LAYER M1 ;
      RECT 12345 15875 12595 16885 ;
    LAYER M1 ;
      RECT 12345 17975 12595 21505 ;
    LAYER M1 ;
      RECT 12345 21755 12595 22765 ;
    LAYER M1 ;
      RECT 12345 23855 12595 27385 ;
    LAYER M1 ;
      RECT 12345 27635 12595 28645 ;
    LAYER M1 ;
      RECT 12345 29735 12595 33265 ;
    LAYER M1 ;
      RECT 12345 33515 12595 34525 ;
    LAYER M1 ;
      RECT 12345 35615 12595 36625 ;
    LAYER M1 ;
      RECT 12775 335 13025 3865 ;
    LAYER M1 ;
      RECT 12775 6215 13025 9745 ;
    LAYER M1 ;
      RECT 12775 12095 13025 15625 ;
    LAYER M1 ;
      RECT 12775 17975 13025 21505 ;
    LAYER M1 ;
      RECT 12775 23855 13025 27385 ;
    LAYER M1 ;
      RECT 12775 29735 13025 33265 ;
    LAYER M1 ;
      RECT 13205 335 13455 3865 ;
    LAYER M1 ;
      RECT 13205 4115 13455 5125 ;
    LAYER M1 ;
      RECT 13205 6215 13455 9745 ;
    LAYER M1 ;
      RECT 13205 9995 13455 11005 ;
    LAYER M1 ;
      RECT 13205 12095 13455 15625 ;
    LAYER M1 ;
      RECT 13205 15875 13455 16885 ;
    LAYER M1 ;
      RECT 13205 17975 13455 21505 ;
    LAYER M1 ;
      RECT 13205 21755 13455 22765 ;
    LAYER M1 ;
      RECT 13205 23855 13455 27385 ;
    LAYER M1 ;
      RECT 13205 27635 13455 28645 ;
    LAYER M1 ;
      RECT 13205 29735 13455 33265 ;
    LAYER M1 ;
      RECT 13205 33515 13455 34525 ;
    LAYER M1 ;
      RECT 13205 35615 13455 36625 ;
    LAYER M1 ;
      RECT 13635 335 13885 3865 ;
    LAYER M1 ;
      RECT 13635 6215 13885 9745 ;
    LAYER M1 ;
      RECT 13635 12095 13885 15625 ;
    LAYER M1 ;
      RECT 13635 17975 13885 21505 ;
    LAYER M1 ;
      RECT 13635 23855 13885 27385 ;
    LAYER M1 ;
      RECT 13635 29735 13885 33265 ;
    LAYER M1 ;
      RECT 14065 335 14315 3865 ;
    LAYER M1 ;
      RECT 14065 4115 14315 5125 ;
    LAYER M1 ;
      RECT 14065 6215 14315 9745 ;
    LAYER M1 ;
      RECT 14065 9995 14315 11005 ;
    LAYER M1 ;
      RECT 14065 12095 14315 15625 ;
    LAYER M1 ;
      RECT 14065 15875 14315 16885 ;
    LAYER M1 ;
      RECT 14065 17975 14315 21505 ;
    LAYER M1 ;
      RECT 14065 21755 14315 22765 ;
    LAYER M1 ;
      RECT 14065 23855 14315 27385 ;
    LAYER M1 ;
      RECT 14065 27635 14315 28645 ;
    LAYER M1 ;
      RECT 14065 29735 14315 33265 ;
    LAYER M1 ;
      RECT 14065 33515 14315 34525 ;
    LAYER M1 ;
      RECT 14065 35615 14315 36625 ;
    LAYER M1 ;
      RECT 14495 335 14745 3865 ;
    LAYER M1 ;
      RECT 14495 6215 14745 9745 ;
    LAYER M1 ;
      RECT 14495 12095 14745 15625 ;
    LAYER M1 ;
      RECT 14495 17975 14745 21505 ;
    LAYER M1 ;
      RECT 14495 23855 14745 27385 ;
    LAYER M1 ;
      RECT 14495 29735 14745 33265 ;
    LAYER M2 ;
      RECT 1120 280 14360 560 ;
    LAYER M2 ;
      RECT 1120 4480 14360 4760 ;
    LAYER M2 ;
      RECT 690 700 14790 980 ;
    LAYER M2 ;
      RECT 1120 6160 14360 6440 ;
    LAYER M2 ;
      RECT 1120 10360 14360 10640 ;
    LAYER M2 ;
      RECT 690 6580 14790 6860 ;
    LAYER M2 ;
      RECT 1120 12040 14360 12320 ;
    LAYER M2 ;
      RECT 1120 16240 14360 16520 ;
    LAYER M2 ;
      RECT 690 12460 14790 12740 ;
    LAYER M2 ;
      RECT 1120 17920 14360 18200 ;
    LAYER M2 ;
      RECT 1120 22120 14360 22400 ;
    LAYER M2 ;
      RECT 690 18340 14790 18620 ;
    LAYER M2 ;
      RECT 1120 23800 14360 24080 ;
    LAYER M2 ;
      RECT 1120 28000 14360 28280 ;
    LAYER M2 ;
      RECT 690 24220 14790 24500 ;
    LAYER M2 ;
      RECT 1120 29680 14360 29960 ;
    LAYER M2 ;
      RECT 1120 33880 14360 34160 ;
    LAYER M2 ;
      RECT 1120 35980 14360 36260 ;
    LAYER M2 ;
      RECT 690 30100 14790 30380 ;
    LAYER V1 ;
      RECT 13245 335 13415 505 ;
    LAYER V1 ;
      RECT 13245 4535 13415 4705 ;
    LAYER V1 ;
      RECT 13245 6215 13415 6385 ;
    LAYER V1 ;
      RECT 13245 10415 13415 10585 ;
    LAYER V1 ;
      RECT 13245 12095 13415 12265 ;
    LAYER V1 ;
      RECT 13245 16295 13415 16465 ;
    LAYER V1 ;
      RECT 13245 17975 13415 18145 ;
    LAYER V1 ;
      RECT 13245 22175 13415 22345 ;
    LAYER V1 ;
      RECT 13245 23855 13415 24025 ;
    LAYER V1 ;
      RECT 13245 28055 13415 28225 ;
    LAYER V1 ;
      RECT 13245 29735 13415 29905 ;
    LAYER V1 ;
      RECT 13245 33935 13415 34105 ;
    LAYER V1 ;
      RECT 13245 36035 13415 36205 ;
    LAYER V1 ;
      RECT 14105 335 14275 505 ;
    LAYER V1 ;
      RECT 14105 4535 14275 4705 ;
    LAYER V1 ;
      RECT 14105 6215 14275 6385 ;
    LAYER V1 ;
      RECT 14105 10415 14275 10585 ;
    LAYER V1 ;
      RECT 14105 12095 14275 12265 ;
    LAYER V1 ;
      RECT 14105 16295 14275 16465 ;
    LAYER V1 ;
      RECT 14105 17975 14275 18145 ;
    LAYER V1 ;
      RECT 14105 22175 14275 22345 ;
    LAYER V1 ;
      RECT 14105 23855 14275 24025 ;
    LAYER V1 ;
      RECT 14105 28055 14275 28225 ;
    LAYER V1 ;
      RECT 14105 29735 14275 29905 ;
    LAYER V1 ;
      RECT 14105 33935 14275 34105 ;
    LAYER V1 ;
      RECT 14105 36035 14275 36205 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 36035 1375 36205 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 29735 2235 29905 ;
    LAYER V1 ;
      RECT 2065 33935 2235 34105 ;
    LAYER V1 ;
      RECT 2065 36035 2235 36205 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12095 3095 12265 ;
    LAYER V1 ;
      RECT 2925 16295 3095 16465 ;
    LAYER V1 ;
      RECT 2925 17975 3095 18145 ;
    LAYER V1 ;
      RECT 2925 22175 3095 22345 ;
    LAYER V1 ;
      RECT 2925 23855 3095 24025 ;
    LAYER V1 ;
      RECT 2925 28055 3095 28225 ;
    LAYER V1 ;
      RECT 2925 29735 3095 29905 ;
    LAYER V1 ;
      RECT 2925 33935 3095 34105 ;
    LAYER V1 ;
      RECT 2925 36035 3095 36205 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12095 3955 12265 ;
    LAYER V1 ;
      RECT 3785 16295 3955 16465 ;
    LAYER V1 ;
      RECT 3785 17975 3955 18145 ;
    LAYER V1 ;
      RECT 3785 22175 3955 22345 ;
    LAYER V1 ;
      RECT 3785 23855 3955 24025 ;
    LAYER V1 ;
      RECT 3785 28055 3955 28225 ;
    LAYER V1 ;
      RECT 3785 29735 3955 29905 ;
    LAYER V1 ;
      RECT 3785 33935 3955 34105 ;
    LAYER V1 ;
      RECT 3785 36035 3955 36205 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12095 4815 12265 ;
    LAYER V1 ;
      RECT 4645 16295 4815 16465 ;
    LAYER V1 ;
      RECT 4645 17975 4815 18145 ;
    LAYER V1 ;
      RECT 4645 22175 4815 22345 ;
    LAYER V1 ;
      RECT 4645 23855 4815 24025 ;
    LAYER V1 ;
      RECT 4645 28055 4815 28225 ;
    LAYER V1 ;
      RECT 4645 29735 4815 29905 ;
    LAYER V1 ;
      RECT 4645 33935 4815 34105 ;
    LAYER V1 ;
      RECT 4645 36035 4815 36205 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12095 5675 12265 ;
    LAYER V1 ;
      RECT 5505 16295 5675 16465 ;
    LAYER V1 ;
      RECT 5505 17975 5675 18145 ;
    LAYER V1 ;
      RECT 5505 22175 5675 22345 ;
    LAYER V1 ;
      RECT 5505 23855 5675 24025 ;
    LAYER V1 ;
      RECT 5505 28055 5675 28225 ;
    LAYER V1 ;
      RECT 5505 29735 5675 29905 ;
    LAYER V1 ;
      RECT 5505 33935 5675 34105 ;
    LAYER V1 ;
      RECT 5505 36035 5675 36205 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6215 6535 6385 ;
    LAYER V1 ;
      RECT 6365 10415 6535 10585 ;
    LAYER V1 ;
      RECT 6365 12095 6535 12265 ;
    LAYER V1 ;
      RECT 6365 16295 6535 16465 ;
    LAYER V1 ;
      RECT 6365 17975 6535 18145 ;
    LAYER V1 ;
      RECT 6365 22175 6535 22345 ;
    LAYER V1 ;
      RECT 6365 23855 6535 24025 ;
    LAYER V1 ;
      RECT 6365 28055 6535 28225 ;
    LAYER V1 ;
      RECT 6365 29735 6535 29905 ;
    LAYER V1 ;
      RECT 6365 33935 6535 34105 ;
    LAYER V1 ;
      RECT 6365 36035 6535 36205 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6215 7395 6385 ;
    LAYER V1 ;
      RECT 7225 10415 7395 10585 ;
    LAYER V1 ;
      RECT 7225 12095 7395 12265 ;
    LAYER V1 ;
      RECT 7225 16295 7395 16465 ;
    LAYER V1 ;
      RECT 7225 17975 7395 18145 ;
    LAYER V1 ;
      RECT 7225 22175 7395 22345 ;
    LAYER V1 ;
      RECT 7225 23855 7395 24025 ;
    LAYER V1 ;
      RECT 7225 28055 7395 28225 ;
    LAYER V1 ;
      RECT 7225 29735 7395 29905 ;
    LAYER V1 ;
      RECT 7225 33935 7395 34105 ;
    LAYER V1 ;
      RECT 7225 36035 7395 36205 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6215 8255 6385 ;
    LAYER V1 ;
      RECT 8085 10415 8255 10585 ;
    LAYER V1 ;
      RECT 8085 12095 8255 12265 ;
    LAYER V1 ;
      RECT 8085 16295 8255 16465 ;
    LAYER V1 ;
      RECT 8085 17975 8255 18145 ;
    LAYER V1 ;
      RECT 8085 22175 8255 22345 ;
    LAYER V1 ;
      RECT 8085 23855 8255 24025 ;
    LAYER V1 ;
      RECT 8085 28055 8255 28225 ;
    LAYER V1 ;
      RECT 8085 29735 8255 29905 ;
    LAYER V1 ;
      RECT 8085 33935 8255 34105 ;
    LAYER V1 ;
      RECT 8085 36035 8255 36205 ;
    LAYER V1 ;
      RECT 8945 335 9115 505 ;
    LAYER V1 ;
      RECT 8945 4535 9115 4705 ;
    LAYER V1 ;
      RECT 8945 6215 9115 6385 ;
    LAYER V1 ;
      RECT 8945 10415 9115 10585 ;
    LAYER V1 ;
      RECT 8945 12095 9115 12265 ;
    LAYER V1 ;
      RECT 8945 16295 9115 16465 ;
    LAYER V1 ;
      RECT 8945 17975 9115 18145 ;
    LAYER V1 ;
      RECT 8945 22175 9115 22345 ;
    LAYER V1 ;
      RECT 8945 23855 9115 24025 ;
    LAYER V1 ;
      RECT 8945 28055 9115 28225 ;
    LAYER V1 ;
      RECT 8945 29735 9115 29905 ;
    LAYER V1 ;
      RECT 8945 33935 9115 34105 ;
    LAYER V1 ;
      RECT 8945 36035 9115 36205 ;
    LAYER V1 ;
      RECT 9805 335 9975 505 ;
    LAYER V1 ;
      RECT 9805 4535 9975 4705 ;
    LAYER V1 ;
      RECT 9805 6215 9975 6385 ;
    LAYER V1 ;
      RECT 9805 10415 9975 10585 ;
    LAYER V1 ;
      RECT 9805 12095 9975 12265 ;
    LAYER V1 ;
      RECT 9805 16295 9975 16465 ;
    LAYER V1 ;
      RECT 9805 17975 9975 18145 ;
    LAYER V1 ;
      RECT 9805 22175 9975 22345 ;
    LAYER V1 ;
      RECT 9805 23855 9975 24025 ;
    LAYER V1 ;
      RECT 9805 28055 9975 28225 ;
    LAYER V1 ;
      RECT 9805 29735 9975 29905 ;
    LAYER V1 ;
      RECT 9805 33935 9975 34105 ;
    LAYER V1 ;
      RECT 9805 36035 9975 36205 ;
    LAYER V1 ;
      RECT 10665 335 10835 505 ;
    LAYER V1 ;
      RECT 10665 4535 10835 4705 ;
    LAYER V1 ;
      RECT 10665 6215 10835 6385 ;
    LAYER V1 ;
      RECT 10665 10415 10835 10585 ;
    LAYER V1 ;
      RECT 10665 12095 10835 12265 ;
    LAYER V1 ;
      RECT 10665 16295 10835 16465 ;
    LAYER V1 ;
      RECT 10665 17975 10835 18145 ;
    LAYER V1 ;
      RECT 10665 22175 10835 22345 ;
    LAYER V1 ;
      RECT 10665 23855 10835 24025 ;
    LAYER V1 ;
      RECT 10665 28055 10835 28225 ;
    LAYER V1 ;
      RECT 10665 29735 10835 29905 ;
    LAYER V1 ;
      RECT 10665 33935 10835 34105 ;
    LAYER V1 ;
      RECT 10665 36035 10835 36205 ;
    LAYER V1 ;
      RECT 11525 335 11695 505 ;
    LAYER V1 ;
      RECT 11525 4535 11695 4705 ;
    LAYER V1 ;
      RECT 11525 6215 11695 6385 ;
    LAYER V1 ;
      RECT 11525 10415 11695 10585 ;
    LAYER V1 ;
      RECT 11525 12095 11695 12265 ;
    LAYER V1 ;
      RECT 11525 16295 11695 16465 ;
    LAYER V1 ;
      RECT 11525 17975 11695 18145 ;
    LAYER V1 ;
      RECT 11525 22175 11695 22345 ;
    LAYER V1 ;
      RECT 11525 23855 11695 24025 ;
    LAYER V1 ;
      RECT 11525 28055 11695 28225 ;
    LAYER V1 ;
      RECT 11525 29735 11695 29905 ;
    LAYER V1 ;
      RECT 11525 33935 11695 34105 ;
    LAYER V1 ;
      RECT 11525 36035 11695 36205 ;
    LAYER V1 ;
      RECT 12385 335 12555 505 ;
    LAYER V1 ;
      RECT 12385 4535 12555 4705 ;
    LAYER V1 ;
      RECT 12385 6215 12555 6385 ;
    LAYER V1 ;
      RECT 12385 10415 12555 10585 ;
    LAYER V1 ;
      RECT 12385 12095 12555 12265 ;
    LAYER V1 ;
      RECT 12385 16295 12555 16465 ;
    LAYER V1 ;
      RECT 12385 17975 12555 18145 ;
    LAYER V1 ;
      RECT 12385 22175 12555 22345 ;
    LAYER V1 ;
      RECT 12385 23855 12555 24025 ;
    LAYER V1 ;
      RECT 12385 28055 12555 28225 ;
    LAYER V1 ;
      RECT 12385 29735 12555 29905 ;
    LAYER V1 ;
      RECT 12385 33935 12555 34105 ;
    LAYER V1 ;
      RECT 12385 36035 12555 36205 ;
    LAYER V1 ;
      RECT 13675 755 13845 925 ;
    LAYER V1 ;
      RECT 13675 6635 13845 6805 ;
    LAYER V1 ;
      RECT 13675 12515 13845 12685 ;
    LAYER V1 ;
      RECT 13675 18395 13845 18565 ;
    LAYER V1 ;
      RECT 13675 24275 13845 24445 ;
    LAYER V1 ;
      RECT 13675 30155 13845 30325 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 14535 755 14705 925 ;
    LAYER V1 ;
      RECT 14535 6635 14705 6805 ;
    LAYER V1 ;
      RECT 14535 12515 14705 12685 ;
    LAYER V1 ;
      RECT 14535 18395 14705 18565 ;
    LAYER V1 ;
      RECT 14535 24275 14705 24445 ;
    LAYER V1 ;
      RECT 14535 30155 14705 30325 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 2495 30155 2665 30325 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 18395 3525 18565 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 3355 30155 3525 30325 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 4215 12515 4385 12685 ;
    LAYER V1 ;
      RECT 4215 18395 4385 18565 ;
    LAYER V1 ;
      RECT 4215 24275 4385 24445 ;
    LAYER V1 ;
      RECT 4215 30155 4385 30325 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 5075 12515 5245 12685 ;
    LAYER V1 ;
      RECT 5075 18395 5245 18565 ;
    LAYER V1 ;
      RECT 5075 24275 5245 24445 ;
    LAYER V1 ;
      RECT 5075 30155 5245 30325 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 5935 6635 6105 6805 ;
    LAYER V1 ;
      RECT 5935 12515 6105 12685 ;
    LAYER V1 ;
      RECT 5935 18395 6105 18565 ;
    LAYER V1 ;
      RECT 5935 24275 6105 24445 ;
    LAYER V1 ;
      RECT 5935 30155 6105 30325 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 6795 12515 6965 12685 ;
    LAYER V1 ;
      RECT 6795 18395 6965 18565 ;
    LAYER V1 ;
      RECT 6795 24275 6965 24445 ;
    LAYER V1 ;
      RECT 6795 30155 6965 30325 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 7655 6635 7825 6805 ;
    LAYER V1 ;
      RECT 7655 12515 7825 12685 ;
    LAYER V1 ;
      RECT 7655 18395 7825 18565 ;
    LAYER V1 ;
      RECT 7655 24275 7825 24445 ;
    LAYER V1 ;
      RECT 7655 30155 7825 30325 ;
    LAYER V1 ;
      RECT 8515 755 8685 925 ;
    LAYER V1 ;
      RECT 8515 6635 8685 6805 ;
    LAYER V1 ;
      RECT 8515 12515 8685 12685 ;
    LAYER V1 ;
      RECT 8515 18395 8685 18565 ;
    LAYER V1 ;
      RECT 8515 24275 8685 24445 ;
    LAYER V1 ;
      RECT 8515 30155 8685 30325 ;
    LAYER V1 ;
      RECT 9375 755 9545 925 ;
    LAYER V1 ;
      RECT 9375 6635 9545 6805 ;
    LAYER V1 ;
      RECT 9375 12515 9545 12685 ;
    LAYER V1 ;
      RECT 9375 18395 9545 18565 ;
    LAYER V1 ;
      RECT 9375 24275 9545 24445 ;
    LAYER V1 ;
      RECT 9375 30155 9545 30325 ;
    LAYER V1 ;
      RECT 10235 755 10405 925 ;
    LAYER V1 ;
      RECT 10235 6635 10405 6805 ;
    LAYER V1 ;
      RECT 10235 12515 10405 12685 ;
    LAYER V1 ;
      RECT 10235 18395 10405 18565 ;
    LAYER V1 ;
      RECT 10235 24275 10405 24445 ;
    LAYER V1 ;
      RECT 10235 30155 10405 30325 ;
    LAYER V1 ;
      RECT 11095 755 11265 925 ;
    LAYER V1 ;
      RECT 11095 6635 11265 6805 ;
    LAYER V1 ;
      RECT 11095 12515 11265 12685 ;
    LAYER V1 ;
      RECT 11095 18395 11265 18565 ;
    LAYER V1 ;
      RECT 11095 24275 11265 24445 ;
    LAYER V1 ;
      RECT 11095 30155 11265 30325 ;
    LAYER V1 ;
      RECT 11955 755 12125 925 ;
    LAYER V1 ;
      RECT 11955 6635 12125 6805 ;
    LAYER V1 ;
      RECT 11955 12515 12125 12685 ;
    LAYER V1 ;
      RECT 11955 18395 12125 18565 ;
    LAYER V1 ;
      RECT 11955 24275 12125 24445 ;
    LAYER V1 ;
      RECT 11955 30155 12125 30325 ;
    LAYER V1 ;
      RECT 12815 755 12985 925 ;
    LAYER V1 ;
      RECT 12815 6635 12985 6805 ;
    LAYER V1 ;
      RECT 12815 12515 12985 12685 ;
    LAYER V1 ;
      RECT 12815 18395 12985 18565 ;
    LAYER V1 ;
      RECT 12815 24275 12985 24445 ;
    LAYER V1 ;
      RECT 12815 30155 12985 30325 ;
    LAYER V2 ;
      RECT 7235 345 7385 495 ;
    LAYER V2 ;
      RECT 7235 6225 7385 6375 ;
    LAYER V2 ;
      RECT 7235 12105 7385 12255 ;
    LAYER V2 ;
      RECT 7235 17985 7385 18135 ;
    LAYER V2 ;
      RECT 7235 23865 7385 24015 ;
    LAYER V2 ;
      RECT 7235 29745 7385 29895 ;
    LAYER V2 ;
      RECT 7665 4545 7815 4695 ;
    LAYER V2 ;
      RECT 7665 10425 7815 10575 ;
    LAYER V2 ;
      RECT 7665 16305 7815 16455 ;
    LAYER V2 ;
      RECT 7665 22185 7815 22335 ;
    LAYER V2 ;
      RECT 7665 28065 7815 28215 ;
    LAYER V2 ;
      RECT 7665 33945 7815 34095 ;
    LAYER V2 ;
      RECT 8095 765 8245 915 ;
    LAYER V2 ;
      RECT 8095 6645 8245 6795 ;
    LAYER V2 ;
      RECT 8095 12525 8245 12675 ;
    LAYER V2 ;
      RECT 8095 18405 8245 18555 ;
    LAYER V2 ;
      RECT 8095 24285 8245 24435 ;
    LAYER V2 ;
      RECT 8095 30165 8245 30315 ;
    LAYER V2 ;
      RECT 8095 36045 8245 36195 ;
  END
END NMOS_S_65192303_X16_Y6
