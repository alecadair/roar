.param w1_2=20.7
.param w3_4=5.00
.param w5_6=90.00
.param w7_8=30.00
.param w9_10=41.4
.param beta=1
.param nf1_2=1
.param nf3_4=1
.param nf5_6=1
.param nf7_8=1
.param nf9_10=1

.param iref_ideal=67.5u
.param iref_post_layout=75u
