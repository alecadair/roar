.param w1_2=11.75
.param w3_4=3.65
.param w5_6=8.06
.param w7_8=25.0
.param w9_10=24.0
.param beta=1
.param nf1_2=1
.param nf3_4=1
.param nf5_6=1
.param nf7_8=1
.param nf9_10=1

.param iref_ideal=65u
.param iref_post_layout=75u
