MACRO NMOS_S_21039285_X1_Y10
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_21039285_X1_Y10 0 0 ;
  SIZE 2580 BY 60480 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720 260 1000 53500 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 4460 1430 57700 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 59800 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 60145 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M2 ;
      RECT 260 280 1460 560 ;
    LAYER M2 ;
      RECT 260 4480 1460 4760 ;
    LAYER M2 ;
      RECT 690 700 1890 980 ;
    LAYER M2 ;
      RECT 260 6160 1460 6440 ;
    LAYER M2 ;
      RECT 260 10360 1460 10640 ;
    LAYER M2 ;
      RECT 690 6580 1890 6860 ;
    LAYER M2 ;
      RECT 260 12040 1460 12320 ;
    LAYER M2 ;
      RECT 260 16240 1460 16520 ;
    LAYER M2 ;
      RECT 690 12460 1890 12740 ;
    LAYER M2 ;
      RECT 260 17920 1460 18200 ;
    LAYER M2 ;
      RECT 260 22120 1460 22400 ;
    LAYER M2 ;
      RECT 690 18340 1890 18620 ;
    LAYER M2 ;
      RECT 260 23800 1460 24080 ;
    LAYER M2 ;
      RECT 260 28000 1460 28280 ;
    LAYER M2 ;
      RECT 690 24220 1890 24500 ;
    LAYER M2 ;
      RECT 260 29680 1460 29960 ;
    LAYER M2 ;
      RECT 260 33880 1460 34160 ;
    LAYER M2 ;
      RECT 690 30100 1890 30380 ;
    LAYER M2 ;
      RECT 260 35560 1460 35840 ;
    LAYER M2 ;
      RECT 260 39760 1460 40040 ;
    LAYER M2 ;
      RECT 690 35980 1890 36260 ;
    LAYER M2 ;
      RECT 260 41440 1460 41720 ;
    LAYER M2 ;
      RECT 260 45640 1460 45920 ;
    LAYER M2 ;
      RECT 690 41860 1890 42140 ;
    LAYER M2 ;
      RECT 260 47320 1460 47600 ;
    LAYER M2 ;
      RECT 260 51520 1460 51800 ;
    LAYER M2 ;
      RECT 690 47740 1890 48020 ;
    LAYER M2 ;
      RECT 260 53200 1460 53480 ;
    LAYER M2 ;
      RECT 260 57400 1460 57680 ;
    LAYER M2 ;
      RECT 690 59500 1890 59780 ;
    LAYER M2 ;
      RECT 690 53620 1890 53900 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53255 1375 53425 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59555 1375 59725 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 775 53675 945 53845 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 1635 53675 1805 53845 ;
    LAYER V2 ;
      RECT 785 345 935 495 ;
    LAYER V2 ;
      RECT 785 6225 935 6375 ;
    LAYER V2 ;
      RECT 785 12105 935 12255 ;
    LAYER V2 ;
      RECT 785 17985 935 18135 ;
    LAYER V2 ;
      RECT 785 23865 935 24015 ;
    LAYER V2 ;
      RECT 785 29745 935 29895 ;
    LAYER V2 ;
      RECT 785 35625 935 35775 ;
    LAYER V2 ;
      RECT 785 41505 935 41655 ;
    LAYER V2 ;
      RECT 785 47385 935 47535 ;
    LAYER V2 ;
      RECT 785 53265 935 53415 ;
    LAYER V2 ;
      RECT 1215 4545 1365 4695 ;
    LAYER V2 ;
      RECT 1215 10425 1365 10575 ;
    LAYER V2 ;
      RECT 1215 16305 1365 16455 ;
    LAYER V2 ;
      RECT 1215 22185 1365 22335 ;
    LAYER V2 ;
      RECT 1215 28065 1365 28215 ;
    LAYER V2 ;
      RECT 1215 33945 1365 34095 ;
    LAYER V2 ;
      RECT 1215 39825 1365 39975 ;
    LAYER V2 ;
      RECT 1215 45705 1365 45855 ;
    LAYER V2 ;
      RECT 1215 51585 1365 51735 ;
    LAYER V2 ;
      RECT 1215 57465 1365 57615 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 6645 1795 6795 ;
    LAYER V2 ;
      RECT 1645 12525 1795 12675 ;
    LAYER V2 ;
      RECT 1645 18405 1795 18555 ;
    LAYER V2 ;
      RECT 1645 24285 1795 24435 ;
    LAYER V2 ;
      RECT 1645 30165 1795 30315 ;
    LAYER V2 ;
      RECT 1645 36045 1795 36195 ;
    LAYER V2 ;
      RECT 1645 41925 1795 42075 ;
    LAYER V2 ;
      RECT 1645 47805 1795 47955 ;
    LAYER V2 ;
      RECT 1645 53685 1795 53835 ;
    LAYER V2 ;
      RECT 1645 59565 1795 59715 ;
  END
END NMOS_S_21039285_X1_Y10
