MACRO NMOS_S_80601593_X5_Y16
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_80601593_X5_Y16 0 0 ;
  SIZE 6020 BY 95760 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 260 2720 88780 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2870 4460 3150 92980 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3300 680 3580 95080 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 62665 ;
    LAYER M1 ;
      RECT 1165 62915 1415 63925 ;
    LAYER M1 ;
      RECT 1165 65015 1415 68545 ;
    LAYER M1 ;
      RECT 1165 68795 1415 69805 ;
    LAYER M1 ;
      RECT 1165 70895 1415 74425 ;
    LAYER M1 ;
      RECT 1165 74675 1415 75685 ;
    LAYER M1 ;
      RECT 1165 76775 1415 80305 ;
    LAYER M1 ;
      RECT 1165 80555 1415 81565 ;
    LAYER M1 ;
      RECT 1165 82655 1415 86185 ;
    LAYER M1 ;
      RECT 1165 86435 1415 87445 ;
    LAYER M1 ;
      RECT 1165 88535 1415 92065 ;
    LAYER M1 ;
      RECT 1165 92315 1415 93325 ;
    LAYER M1 ;
      RECT 1165 94415 1415 95425 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 735 59135 985 62665 ;
    LAYER M1 ;
      RECT 735 65015 985 68545 ;
    LAYER M1 ;
      RECT 735 70895 985 74425 ;
    LAYER M1 ;
      RECT 735 76775 985 80305 ;
    LAYER M1 ;
      RECT 735 82655 985 86185 ;
    LAYER M1 ;
      RECT 735 88535 985 92065 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M1 ;
      RECT 1595 59135 1845 62665 ;
    LAYER M1 ;
      RECT 1595 65015 1845 68545 ;
    LAYER M1 ;
      RECT 1595 70895 1845 74425 ;
    LAYER M1 ;
      RECT 1595 76775 1845 80305 ;
    LAYER M1 ;
      RECT 1595 82655 1845 86185 ;
    LAYER M1 ;
      RECT 1595 88535 1845 92065 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 33265 ;
    LAYER M1 ;
      RECT 2025 33515 2275 34525 ;
    LAYER M1 ;
      RECT 2025 35615 2275 39145 ;
    LAYER M1 ;
      RECT 2025 39395 2275 40405 ;
    LAYER M1 ;
      RECT 2025 41495 2275 45025 ;
    LAYER M1 ;
      RECT 2025 45275 2275 46285 ;
    LAYER M1 ;
      RECT 2025 47375 2275 50905 ;
    LAYER M1 ;
      RECT 2025 51155 2275 52165 ;
    LAYER M1 ;
      RECT 2025 53255 2275 56785 ;
    LAYER M1 ;
      RECT 2025 57035 2275 58045 ;
    LAYER M1 ;
      RECT 2025 59135 2275 62665 ;
    LAYER M1 ;
      RECT 2025 62915 2275 63925 ;
    LAYER M1 ;
      RECT 2025 65015 2275 68545 ;
    LAYER M1 ;
      RECT 2025 68795 2275 69805 ;
    LAYER M1 ;
      RECT 2025 70895 2275 74425 ;
    LAYER M1 ;
      RECT 2025 74675 2275 75685 ;
    LAYER M1 ;
      RECT 2025 76775 2275 80305 ;
    LAYER M1 ;
      RECT 2025 80555 2275 81565 ;
    LAYER M1 ;
      RECT 2025 82655 2275 86185 ;
    LAYER M1 ;
      RECT 2025 86435 2275 87445 ;
    LAYER M1 ;
      RECT 2025 88535 2275 92065 ;
    LAYER M1 ;
      RECT 2025 92315 2275 93325 ;
    LAYER M1 ;
      RECT 2025 94415 2275 95425 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2455 35615 2705 39145 ;
    LAYER M1 ;
      RECT 2455 41495 2705 45025 ;
    LAYER M1 ;
      RECT 2455 47375 2705 50905 ;
    LAYER M1 ;
      RECT 2455 53255 2705 56785 ;
    LAYER M1 ;
      RECT 2455 59135 2705 62665 ;
    LAYER M1 ;
      RECT 2455 65015 2705 68545 ;
    LAYER M1 ;
      RECT 2455 70895 2705 74425 ;
    LAYER M1 ;
      RECT 2455 76775 2705 80305 ;
    LAYER M1 ;
      RECT 2455 82655 2705 86185 ;
    LAYER M1 ;
      RECT 2455 88535 2705 92065 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 15625 ;
    LAYER M1 ;
      RECT 2885 15875 3135 16885 ;
    LAYER M1 ;
      RECT 2885 17975 3135 21505 ;
    LAYER M1 ;
      RECT 2885 21755 3135 22765 ;
    LAYER M1 ;
      RECT 2885 23855 3135 27385 ;
    LAYER M1 ;
      RECT 2885 27635 3135 28645 ;
    LAYER M1 ;
      RECT 2885 29735 3135 33265 ;
    LAYER M1 ;
      RECT 2885 33515 3135 34525 ;
    LAYER M1 ;
      RECT 2885 35615 3135 39145 ;
    LAYER M1 ;
      RECT 2885 39395 3135 40405 ;
    LAYER M1 ;
      RECT 2885 41495 3135 45025 ;
    LAYER M1 ;
      RECT 2885 45275 3135 46285 ;
    LAYER M1 ;
      RECT 2885 47375 3135 50905 ;
    LAYER M1 ;
      RECT 2885 51155 3135 52165 ;
    LAYER M1 ;
      RECT 2885 53255 3135 56785 ;
    LAYER M1 ;
      RECT 2885 57035 3135 58045 ;
    LAYER M1 ;
      RECT 2885 59135 3135 62665 ;
    LAYER M1 ;
      RECT 2885 62915 3135 63925 ;
    LAYER M1 ;
      RECT 2885 65015 3135 68545 ;
    LAYER M1 ;
      RECT 2885 68795 3135 69805 ;
    LAYER M1 ;
      RECT 2885 70895 3135 74425 ;
    LAYER M1 ;
      RECT 2885 74675 3135 75685 ;
    LAYER M1 ;
      RECT 2885 76775 3135 80305 ;
    LAYER M1 ;
      RECT 2885 80555 3135 81565 ;
    LAYER M1 ;
      RECT 2885 82655 3135 86185 ;
    LAYER M1 ;
      RECT 2885 86435 3135 87445 ;
    LAYER M1 ;
      RECT 2885 88535 3135 92065 ;
    LAYER M1 ;
      RECT 2885 92315 3135 93325 ;
    LAYER M1 ;
      RECT 2885 94415 3135 95425 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 23855 3565 27385 ;
    LAYER M1 ;
      RECT 3315 29735 3565 33265 ;
    LAYER M1 ;
      RECT 3315 35615 3565 39145 ;
    LAYER M1 ;
      RECT 3315 41495 3565 45025 ;
    LAYER M1 ;
      RECT 3315 47375 3565 50905 ;
    LAYER M1 ;
      RECT 3315 53255 3565 56785 ;
    LAYER M1 ;
      RECT 3315 59135 3565 62665 ;
    LAYER M1 ;
      RECT 3315 65015 3565 68545 ;
    LAYER M1 ;
      RECT 3315 70895 3565 74425 ;
    LAYER M1 ;
      RECT 3315 76775 3565 80305 ;
    LAYER M1 ;
      RECT 3315 82655 3565 86185 ;
    LAYER M1 ;
      RECT 3315 88535 3565 92065 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 15625 ;
    LAYER M1 ;
      RECT 3745 15875 3995 16885 ;
    LAYER M1 ;
      RECT 3745 17975 3995 21505 ;
    LAYER M1 ;
      RECT 3745 21755 3995 22765 ;
    LAYER M1 ;
      RECT 3745 23855 3995 27385 ;
    LAYER M1 ;
      RECT 3745 27635 3995 28645 ;
    LAYER M1 ;
      RECT 3745 29735 3995 33265 ;
    LAYER M1 ;
      RECT 3745 33515 3995 34525 ;
    LAYER M1 ;
      RECT 3745 35615 3995 39145 ;
    LAYER M1 ;
      RECT 3745 39395 3995 40405 ;
    LAYER M1 ;
      RECT 3745 41495 3995 45025 ;
    LAYER M1 ;
      RECT 3745 45275 3995 46285 ;
    LAYER M1 ;
      RECT 3745 47375 3995 50905 ;
    LAYER M1 ;
      RECT 3745 51155 3995 52165 ;
    LAYER M1 ;
      RECT 3745 53255 3995 56785 ;
    LAYER M1 ;
      RECT 3745 57035 3995 58045 ;
    LAYER M1 ;
      RECT 3745 59135 3995 62665 ;
    LAYER M1 ;
      RECT 3745 62915 3995 63925 ;
    LAYER M1 ;
      RECT 3745 65015 3995 68545 ;
    LAYER M1 ;
      RECT 3745 68795 3995 69805 ;
    LAYER M1 ;
      RECT 3745 70895 3995 74425 ;
    LAYER M1 ;
      RECT 3745 74675 3995 75685 ;
    LAYER M1 ;
      RECT 3745 76775 3995 80305 ;
    LAYER M1 ;
      RECT 3745 80555 3995 81565 ;
    LAYER M1 ;
      RECT 3745 82655 3995 86185 ;
    LAYER M1 ;
      RECT 3745 86435 3995 87445 ;
    LAYER M1 ;
      RECT 3745 88535 3995 92065 ;
    LAYER M1 ;
      RECT 3745 92315 3995 93325 ;
    LAYER M1 ;
      RECT 3745 94415 3995 95425 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4175 17975 4425 21505 ;
    LAYER M1 ;
      RECT 4175 23855 4425 27385 ;
    LAYER M1 ;
      RECT 4175 29735 4425 33265 ;
    LAYER M1 ;
      RECT 4175 35615 4425 39145 ;
    LAYER M1 ;
      RECT 4175 41495 4425 45025 ;
    LAYER M1 ;
      RECT 4175 47375 4425 50905 ;
    LAYER M1 ;
      RECT 4175 53255 4425 56785 ;
    LAYER M1 ;
      RECT 4175 59135 4425 62665 ;
    LAYER M1 ;
      RECT 4175 65015 4425 68545 ;
    LAYER M1 ;
      RECT 4175 70895 4425 74425 ;
    LAYER M1 ;
      RECT 4175 76775 4425 80305 ;
    LAYER M1 ;
      RECT 4175 82655 4425 86185 ;
    LAYER M1 ;
      RECT 4175 88535 4425 92065 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 15625 ;
    LAYER M1 ;
      RECT 4605 15875 4855 16885 ;
    LAYER M1 ;
      RECT 4605 17975 4855 21505 ;
    LAYER M1 ;
      RECT 4605 21755 4855 22765 ;
    LAYER M1 ;
      RECT 4605 23855 4855 27385 ;
    LAYER M1 ;
      RECT 4605 27635 4855 28645 ;
    LAYER M1 ;
      RECT 4605 29735 4855 33265 ;
    LAYER M1 ;
      RECT 4605 33515 4855 34525 ;
    LAYER M1 ;
      RECT 4605 35615 4855 39145 ;
    LAYER M1 ;
      RECT 4605 39395 4855 40405 ;
    LAYER M1 ;
      RECT 4605 41495 4855 45025 ;
    LAYER M1 ;
      RECT 4605 45275 4855 46285 ;
    LAYER M1 ;
      RECT 4605 47375 4855 50905 ;
    LAYER M1 ;
      RECT 4605 51155 4855 52165 ;
    LAYER M1 ;
      RECT 4605 53255 4855 56785 ;
    LAYER M1 ;
      RECT 4605 57035 4855 58045 ;
    LAYER M1 ;
      RECT 4605 59135 4855 62665 ;
    LAYER M1 ;
      RECT 4605 62915 4855 63925 ;
    LAYER M1 ;
      RECT 4605 65015 4855 68545 ;
    LAYER M1 ;
      RECT 4605 68795 4855 69805 ;
    LAYER M1 ;
      RECT 4605 70895 4855 74425 ;
    LAYER M1 ;
      RECT 4605 74675 4855 75685 ;
    LAYER M1 ;
      RECT 4605 76775 4855 80305 ;
    LAYER M1 ;
      RECT 4605 80555 4855 81565 ;
    LAYER M1 ;
      RECT 4605 82655 4855 86185 ;
    LAYER M1 ;
      RECT 4605 86435 4855 87445 ;
    LAYER M1 ;
      RECT 4605 88535 4855 92065 ;
    LAYER M1 ;
      RECT 4605 92315 4855 93325 ;
    LAYER M1 ;
      RECT 4605 94415 4855 95425 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5035 12095 5285 15625 ;
    LAYER M1 ;
      RECT 5035 17975 5285 21505 ;
    LAYER M1 ;
      RECT 5035 23855 5285 27385 ;
    LAYER M1 ;
      RECT 5035 29735 5285 33265 ;
    LAYER M1 ;
      RECT 5035 35615 5285 39145 ;
    LAYER M1 ;
      RECT 5035 41495 5285 45025 ;
    LAYER M1 ;
      RECT 5035 47375 5285 50905 ;
    LAYER M1 ;
      RECT 5035 53255 5285 56785 ;
    LAYER M1 ;
      RECT 5035 59135 5285 62665 ;
    LAYER M1 ;
      RECT 5035 65015 5285 68545 ;
    LAYER M1 ;
      RECT 5035 70895 5285 74425 ;
    LAYER M1 ;
      RECT 5035 76775 5285 80305 ;
    LAYER M1 ;
      RECT 5035 82655 5285 86185 ;
    LAYER M1 ;
      RECT 5035 88535 5285 92065 ;
    LAYER M2 ;
      RECT 1120 280 4900 560 ;
    LAYER M2 ;
      RECT 1120 4480 4900 4760 ;
    LAYER M2 ;
      RECT 690 700 5330 980 ;
    LAYER M2 ;
      RECT 1120 6160 4900 6440 ;
    LAYER M2 ;
      RECT 1120 10360 4900 10640 ;
    LAYER M2 ;
      RECT 690 6580 5330 6860 ;
    LAYER M2 ;
      RECT 1120 12040 4900 12320 ;
    LAYER M2 ;
      RECT 1120 16240 4900 16520 ;
    LAYER M2 ;
      RECT 690 12460 5330 12740 ;
    LAYER M2 ;
      RECT 1120 17920 4900 18200 ;
    LAYER M2 ;
      RECT 1120 22120 4900 22400 ;
    LAYER M2 ;
      RECT 690 18340 5330 18620 ;
    LAYER M2 ;
      RECT 1120 23800 4900 24080 ;
    LAYER M2 ;
      RECT 1120 28000 4900 28280 ;
    LAYER M2 ;
      RECT 690 24220 5330 24500 ;
    LAYER M2 ;
      RECT 1120 29680 4900 29960 ;
    LAYER M2 ;
      RECT 1120 33880 4900 34160 ;
    LAYER M2 ;
      RECT 690 30100 5330 30380 ;
    LAYER M2 ;
      RECT 1120 35560 4900 35840 ;
    LAYER M2 ;
      RECT 1120 39760 4900 40040 ;
    LAYER M2 ;
      RECT 690 35980 5330 36260 ;
    LAYER M2 ;
      RECT 1120 41440 4900 41720 ;
    LAYER M2 ;
      RECT 1120 45640 4900 45920 ;
    LAYER M2 ;
      RECT 690 41860 5330 42140 ;
    LAYER M2 ;
      RECT 1120 47320 4900 47600 ;
    LAYER M2 ;
      RECT 1120 51520 4900 51800 ;
    LAYER M2 ;
      RECT 690 47740 5330 48020 ;
    LAYER M2 ;
      RECT 1120 53200 4900 53480 ;
    LAYER M2 ;
      RECT 1120 57400 4900 57680 ;
    LAYER M2 ;
      RECT 690 53620 5330 53900 ;
    LAYER M2 ;
      RECT 1120 59080 4900 59360 ;
    LAYER M2 ;
      RECT 1120 63280 4900 63560 ;
    LAYER M2 ;
      RECT 690 59500 5330 59780 ;
    LAYER M2 ;
      RECT 1120 64960 4900 65240 ;
    LAYER M2 ;
      RECT 1120 69160 4900 69440 ;
    LAYER M2 ;
      RECT 690 65380 5330 65660 ;
    LAYER M2 ;
      RECT 1120 70840 4900 71120 ;
    LAYER M2 ;
      RECT 1120 75040 4900 75320 ;
    LAYER M2 ;
      RECT 690 71260 5330 71540 ;
    LAYER M2 ;
      RECT 1120 76720 4900 77000 ;
    LAYER M2 ;
      RECT 1120 80920 4900 81200 ;
    LAYER M2 ;
      RECT 690 77140 5330 77420 ;
    LAYER M2 ;
      RECT 1120 82600 4900 82880 ;
    LAYER M2 ;
      RECT 1120 86800 4900 87080 ;
    LAYER M2 ;
      RECT 690 83020 5330 83300 ;
    LAYER M2 ;
      RECT 1120 88480 4900 88760 ;
    LAYER M2 ;
      RECT 1120 92680 4900 92960 ;
    LAYER M2 ;
      RECT 1120 94780 4900 95060 ;
    LAYER M2 ;
      RECT 690 88900 5330 89180 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53255 1375 53425 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59135 1375 59305 ;
    LAYER V1 ;
      RECT 1205 63335 1375 63505 ;
    LAYER V1 ;
      RECT 1205 65015 1375 65185 ;
    LAYER V1 ;
      RECT 1205 69215 1375 69385 ;
    LAYER V1 ;
      RECT 1205 70895 1375 71065 ;
    LAYER V1 ;
      RECT 1205 75095 1375 75265 ;
    LAYER V1 ;
      RECT 1205 76775 1375 76945 ;
    LAYER V1 ;
      RECT 1205 80975 1375 81145 ;
    LAYER V1 ;
      RECT 1205 82655 1375 82825 ;
    LAYER V1 ;
      RECT 1205 86855 1375 87025 ;
    LAYER V1 ;
      RECT 1205 88535 1375 88705 ;
    LAYER V1 ;
      RECT 1205 92735 1375 92905 ;
    LAYER V1 ;
      RECT 1205 94835 1375 95005 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 29735 2235 29905 ;
    LAYER V1 ;
      RECT 2065 33935 2235 34105 ;
    LAYER V1 ;
      RECT 2065 35615 2235 35785 ;
    LAYER V1 ;
      RECT 2065 39815 2235 39985 ;
    LAYER V1 ;
      RECT 2065 41495 2235 41665 ;
    LAYER V1 ;
      RECT 2065 45695 2235 45865 ;
    LAYER V1 ;
      RECT 2065 47375 2235 47545 ;
    LAYER V1 ;
      RECT 2065 51575 2235 51745 ;
    LAYER V1 ;
      RECT 2065 53255 2235 53425 ;
    LAYER V1 ;
      RECT 2065 57455 2235 57625 ;
    LAYER V1 ;
      RECT 2065 59135 2235 59305 ;
    LAYER V1 ;
      RECT 2065 63335 2235 63505 ;
    LAYER V1 ;
      RECT 2065 65015 2235 65185 ;
    LAYER V1 ;
      RECT 2065 69215 2235 69385 ;
    LAYER V1 ;
      RECT 2065 70895 2235 71065 ;
    LAYER V1 ;
      RECT 2065 75095 2235 75265 ;
    LAYER V1 ;
      RECT 2065 76775 2235 76945 ;
    LAYER V1 ;
      RECT 2065 80975 2235 81145 ;
    LAYER V1 ;
      RECT 2065 82655 2235 82825 ;
    LAYER V1 ;
      RECT 2065 86855 2235 87025 ;
    LAYER V1 ;
      RECT 2065 88535 2235 88705 ;
    LAYER V1 ;
      RECT 2065 92735 2235 92905 ;
    LAYER V1 ;
      RECT 2065 94835 2235 95005 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12095 3095 12265 ;
    LAYER V1 ;
      RECT 2925 16295 3095 16465 ;
    LAYER V1 ;
      RECT 2925 17975 3095 18145 ;
    LAYER V1 ;
      RECT 2925 22175 3095 22345 ;
    LAYER V1 ;
      RECT 2925 23855 3095 24025 ;
    LAYER V1 ;
      RECT 2925 28055 3095 28225 ;
    LAYER V1 ;
      RECT 2925 29735 3095 29905 ;
    LAYER V1 ;
      RECT 2925 33935 3095 34105 ;
    LAYER V1 ;
      RECT 2925 35615 3095 35785 ;
    LAYER V1 ;
      RECT 2925 39815 3095 39985 ;
    LAYER V1 ;
      RECT 2925 41495 3095 41665 ;
    LAYER V1 ;
      RECT 2925 45695 3095 45865 ;
    LAYER V1 ;
      RECT 2925 47375 3095 47545 ;
    LAYER V1 ;
      RECT 2925 51575 3095 51745 ;
    LAYER V1 ;
      RECT 2925 53255 3095 53425 ;
    LAYER V1 ;
      RECT 2925 57455 3095 57625 ;
    LAYER V1 ;
      RECT 2925 59135 3095 59305 ;
    LAYER V1 ;
      RECT 2925 63335 3095 63505 ;
    LAYER V1 ;
      RECT 2925 65015 3095 65185 ;
    LAYER V1 ;
      RECT 2925 69215 3095 69385 ;
    LAYER V1 ;
      RECT 2925 70895 3095 71065 ;
    LAYER V1 ;
      RECT 2925 75095 3095 75265 ;
    LAYER V1 ;
      RECT 2925 76775 3095 76945 ;
    LAYER V1 ;
      RECT 2925 80975 3095 81145 ;
    LAYER V1 ;
      RECT 2925 82655 3095 82825 ;
    LAYER V1 ;
      RECT 2925 86855 3095 87025 ;
    LAYER V1 ;
      RECT 2925 88535 3095 88705 ;
    LAYER V1 ;
      RECT 2925 92735 3095 92905 ;
    LAYER V1 ;
      RECT 2925 94835 3095 95005 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12095 3955 12265 ;
    LAYER V1 ;
      RECT 3785 16295 3955 16465 ;
    LAYER V1 ;
      RECT 3785 17975 3955 18145 ;
    LAYER V1 ;
      RECT 3785 22175 3955 22345 ;
    LAYER V1 ;
      RECT 3785 23855 3955 24025 ;
    LAYER V1 ;
      RECT 3785 28055 3955 28225 ;
    LAYER V1 ;
      RECT 3785 29735 3955 29905 ;
    LAYER V1 ;
      RECT 3785 33935 3955 34105 ;
    LAYER V1 ;
      RECT 3785 35615 3955 35785 ;
    LAYER V1 ;
      RECT 3785 39815 3955 39985 ;
    LAYER V1 ;
      RECT 3785 41495 3955 41665 ;
    LAYER V1 ;
      RECT 3785 45695 3955 45865 ;
    LAYER V1 ;
      RECT 3785 47375 3955 47545 ;
    LAYER V1 ;
      RECT 3785 51575 3955 51745 ;
    LAYER V1 ;
      RECT 3785 53255 3955 53425 ;
    LAYER V1 ;
      RECT 3785 57455 3955 57625 ;
    LAYER V1 ;
      RECT 3785 59135 3955 59305 ;
    LAYER V1 ;
      RECT 3785 63335 3955 63505 ;
    LAYER V1 ;
      RECT 3785 65015 3955 65185 ;
    LAYER V1 ;
      RECT 3785 69215 3955 69385 ;
    LAYER V1 ;
      RECT 3785 70895 3955 71065 ;
    LAYER V1 ;
      RECT 3785 75095 3955 75265 ;
    LAYER V1 ;
      RECT 3785 76775 3955 76945 ;
    LAYER V1 ;
      RECT 3785 80975 3955 81145 ;
    LAYER V1 ;
      RECT 3785 82655 3955 82825 ;
    LAYER V1 ;
      RECT 3785 86855 3955 87025 ;
    LAYER V1 ;
      RECT 3785 88535 3955 88705 ;
    LAYER V1 ;
      RECT 3785 92735 3955 92905 ;
    LAYER V1 ;
      RECT 3785 94835 3955 95005 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12095 4815 12265 ;
    LAYER V1 ;
      RECT 4645 16295 4815 16465 ;
    LAYER V1 ;
      RECT 4645 17975 4815 18145 ;
    LAYER V1 ;
      RECT 4645 22175 4815 22345 ;
    LAYER V1 ;
      RECT 4645 23855 4815 24025 ;
    LAYER V1 ;
      RECT 4645 28055 4815 28225 ;
    LAYER V1 ;
      RECT 4645 29735 4815 29905 ;
    LAYER V1 ;
      RECT 4645 33935 4815 34105 ;
    LAYER V1 ;
      RECT 4645 35615 4815 35785 ;
    LAYER V1 ;
      RECT 4645 39815 4815 39985 ;
    LAYER V1 ;
      RECT 4645 41495 4815 41665 ;
    LAYER V1 ;
      RECT 4645 45695 4815 45865 ;
    LAYER V1 ;
      RECT 4645 47375 4815 47545 ;
    LAYER V1 ;
      RECT 4645 51575 4815 51745 ;
    LAYER V1 ;
      RECT 4645 53255 4815 53425 ;
    LAYER V1 ;
      RECT 4645 57455 4815 57625 ;
    LAYER V1 ;
      RECT 4645 59135 4815 59305 ;
    LAYER V1 ;
      RECT 4645 63335 4815 63505 ;
    LAYER V1 ;
      RECT 4645 65015 4815 65185 ;
    LAYER V1 ;
      RECT 4645 69215 4815 69385 ;
    LAYER V1 ;
      RECT 4645 70895 4815 71065 ;
    LAYER V1 ;
      RECT 4645 75095 4815 75265 ;
    LAYER V1 ;
      RECT 4645 76775 4815 76945 ;
    LAYER V1 ;
      RECT 4645 80975 4815 81145 ;
    LAYER V1 ;
      RECT 4645 82655 4815 82825 ;
    LAYER V1 ;
      RECT 4645 86855 4815 87025 ;
    LAYER V1 ;
      RECT 4645 88535 4815 88705 ;
    LAYER V1 ;
      RECT 4645 92735 4815 92905 ;
    LAYER V1 ;
      RECT 4645 94835 4815 95005 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 775 53675 945 53845 ;
    LAYER V1 ;
      RECT 775 59555 945 59725 ;
    LAYER V1 ;
      RECT 775 65435 945 65605 ;
    LAYER V1 ;
      RECT 775 71315 945 71485 ;
    LAYER V1 ;
      RECT 775 77195 945 77365 ;
    LAYER V1 ;
      RECT 775 83075 945 83245 ;
    LAYER V1 ;
      RECT 775 88955 945 89125 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 1635 53675 1805 53845 ;
    LAYER V1 ;
      RECT 1635 59555 1805 59725 ;
    LAYER V1 ;
      RECT 1635 65435 1805 65605 ;
    LAYER V1 ;
      RECT 1635 71315 1805 71485 ;
    LAYER V1 ;
      RECT 1635 77195 1805 77365 ;
    LAYER V1 ;
      RECT 1635 83075 1805 83245 ;
    LAYER V1 ;
      RECT 1635 88955 1805 89125 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 2495 30155 2665 30325 ;
    LAYER V1 ;
      RECT 2495 36035 2665 36205 ;
    LAYER V1 ;
      RECT 2495 41915 2665 42085 ;
    LAYER V1 ;
      RECT 2495 47795 2665 47965 ;
    LAYER V1 ;
      RECT 2495 53675 2665 53845 ;
    LAYER V1 ;
      RECT 2495 59555 2665 59725 ;
    LAYER V1 ;
      RECT 2495 65435 2665 65605 ;
    LAYER V1 ;
      RECT 2495 71315 2665 71485 ;
    LAYER V1 ;
      RECT 2495 77195 2665 77365 ;
    LAYER V1 ;
      RECT 2495 83075 2665 83245 ;
    LAYER V1 ;
      RECT 2495 88955 2665 89125 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 18395 3525 18565 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 3355 30155 3525 30325 ;
    LAYER V1 ;
      RECT 3355 36035 3525 36205 ;
    LAYER V1 ;
      RECT 3355 41915 3525 42085 ;
    LAYER V1 ;
      RECT 3355 47795 3525 47965 ;
    LAYER V1 ;
      RECT 3355 53675 3525 53845 ;
    LAYER V1 ;
      RECT 3355 59555 3525 59725 ;
    LAYER V1 ;
      RECT 3355 65435 3525 65605 ;
    LAYER V1 ;
      RECT 3355 71315 3525 71485 ;
    LAYER V1 ;
      RECT 3355 77195 3525 77365 ;
    LAYER V1 ;
      RECT 3355 83075 3525 83245 ;
    LAYER V1 ;
      RECT 3355 88955 3525 89125 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 4215 12515 4385 12685 ;
    LAYER V1 ;
      RECT 4215 18395 4385 18565 ;
    LAYER V1 ;
      RECT 4215 24275 4385 24445 ;
    LAYER V1 ;
      RECT 4215 30155 4385 30325 ;
    LAYER V1 ;
      RECT 4215 36035 4385 36205 ;
    LAYER V1 ;
      RECT 4215 41915 4385 42085 ;
    LAYER V1 ;
      RECT 4215 47795 4385 47965 ;
    LAYER V1 ;
      RECT 4215 53675 4385 53845 ;
    LAYER V1 ;
      RECT 4215 59555 4385 59725 ;
    LAYER V1 ;
      RECT 4215 65435 4385 65605 ;
    LAYER V1 ;
      RECT 4215 71315 4385 71485 ;
    LAYER V1 ;
      RECT 4215 77195 4385 77365 ;
    LAYER V1 ;
      RECT 4215 83075 4385 83245 ;
    LAYER V1 ;
      RECT 4215 88955 4385 89125 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 5075 12515 5245 12685 ;
    LAYER V1 ;
      RECT 5075 18395 5245 18565 ;
    LAYER V1 ;
      RECT 5075 24275 5245 24445 ;
    LAYER V1 ;
      RECT 5075 30155 5245 30325 ;
    LAYER V1 ;
      RECT 5075 36035 5245 36205 ;
    LAYER V1 ;
      RECT 5075 41915 5245 42085 ;
    LAYER V1 ;
      RECT 5075 47795 5245 47965 ;
    LAYER V1 ;
      RECT 5075 53675 5245 53845 ;
    LAYER V1 ;
      RECT 5075 59555 5245 59725 ;
    LAYER V1 ;
      RECT 5075 65435 5245 65605 ;
    LAYER V1 ;
      RECT 5075 71315 5245 71485 ;
    LAYER V1 ;
      RECT 5075 77195 5245 77365 ;
    LAYER V1 ;
      RECT 5075 83075 5245 83245 ;
    LAYER V1 ;
      RECT 5075 88955 5245 89125 ;
    LAYER V2 ;
      RECT 2505 345 2655 495 ;
    LAYER V2 ;
      RECT 2505 6225 2655 6375 ;
    LAYER V2 ;
      RECT 2505 12105 2655 12255 ;
    LAYER V2 ;
      RECT 2505 17985 2655 18135 ;
    LAYER V2 ;
      RECT 2505 23865 2655 24015 ;
    LAYER V2 ;
      RECT 2505 29745 2655 29895 ;
    LAYER V2 ;
      RECT 2505 35625 2655 35775 ;
    LAYER V2 ;
      RECT 2505 41505 2655 41655 ;
    LAYER V2 ;
      RECT 2505 47385 2655 47535 ;
    LAYER V2 ;
      RECT 2505 53265 2655 53415 ;
    LAYER V2 ;
      RECT 2505 59145 2655 59295 ;
    LAYER V2 ;
      RECT 2505 65025 2655 65175 ;
    LAYER V2 ;
      RECT 2505 70905 2655 71055 ;
    LAYER V2 ;
      RECT 2505 76785 2655 76935 ;
    LAYER V2 ;
      RECT 2505 82665 2655 82815 ;
    LAYER V2 ;
      RECT 2505 88545 2655 88695 ;
    LAYER V2 ;
      RECT 2935 4545 3085 4695 ;
    LAYER V2 ;
      RECT 2935 10425 3085 10575 ;
    LAYER V2 ;
      RECT 2935 16305 3085 16455 ;
    LAYER V2 ;
      RECT 2935 22185 3085 22335 ;
    LAYER V2 ;
      RECT 2935 28065 3085 28215 ;
    LAYER V2 ;
      RECT 2935 33945 3085 34095 ;
    LAYER V2 ;
      RECT 2935 39825 3085 39975 ;
    LAYER V2 ;
      RECT 2935 45705 3085 45855 ;
    LAYER V2 ;
      RECT 2935 51585 3085 51735 ;
    LAYER V2 ;
      RECT 2935 57465 3085 57615 ;
    LAYER V2 ;
      RECT 2935 63345 3085 63495 ;
    LAYER V2 ;
      RECT 2935 69225 3085 69375 ;
    LAYER V2 ;
      RECT 2935 75105 3085 75255 ;
    LAYER V2 ;
      RECT 2935 80985 3085 81135 ;
    LAYER V2 ;
      RECT 2935 86865 3085 87015 ;
    LAYER V2 ;
      RECT 2935 92745 3085 92895 ;
    LAYER V2 ;
      RECT 3365 765 3515 915 ;
    LAYER V2 ;
      RECT 3365 6645 3515 6795 ;
    LAYER V2 ;
      RECT 3365 12525 3515 12675 ;
    LAYER V2 ;
      RECT 3365 18405 3515 18555 ;
    LAYER V2 ;
      RECT 3365 24285 3515 24435 ;
    LAYER V2 ;
      RECT 3365 30165 3515 30315 ;
    LAYER V2 ;
      RECT 3365 36045 3515 36195 ;
    LAYER V2 ;
      RECT 3365 41925 3515 42075 ;
    LAYER V2 ;
      RECT 3365 47805 3515 47955 ;
    LAYER V2 ;
      RECT 3365 53685 3515 53835 ;
    LAYER V2 ;
      RECT 3365 59565 3515 59715 ;
    LAYER V2 ;
      RECT 3365 65445 3515 65595 ;
    LAYER V2 ;
      RECT 3365 71325 3515 71475 ;
    LAYER V2 ;
      RECT 3365 77205 3515 77355 ;
    LAYER V2 ;
      RECT 3365 83085 3515 83235 ;
    LAYER V2 ;
      RECT 3365 88965 3515 89115 ;
    LAYER V2 ;
      RECT 3365 94845 3515 94995 ;
  END
END NMOS_S_80601593_X5_Y16
