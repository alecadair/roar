MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 38.83 BY 46.79 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 13.62 2.78 13.9 7.3 ;
      LAYER M2 ;
        RECT 20.04 2.8 28.12 3.08 ;
      LAYER M3 ;
        RECT 13.62 3.175 13.9 3.545 ;
      LAYER M2 ;
        RECT 13.76 3.22 18.92 3.5 ;
      LAYER M1 ;
        RECT 18.795 2.94 19.045 3.36 ;
      LAYER M2 ;
        RECT 18.92 2.8 20.21 3.08 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 7.17 14.54 7.45 20.74 ;
      LAYER M3 ;
        RECT 8.89 21.26 9.17 39.22 ;
      LAYER M3 ;
        RECT 7.17 20.58 7.45 21.42 ;
      LAYER M4 ;
        RECT 7.31 21.02 9.03 21.82 ;
      LAYER M3 ;
        RECT 8.89 21.235 9.17 21.605 ;
    END
  END VOUT
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 21.79 12.02 22.07 18.22 ;
    END
  END VINN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 15.77 12.02 16.05 18.22 ;
    END
  END VINP
  OBS 
  LAYER M3 ;
        RECT 9.32 25.46 9.6 43.42 ;
  LAYER M3 ;
        RECT 28.24 21.26 28.52 43.42 ;
  LAYER M3 ;
        RECT 30.39 14.54 30.67 20.74 ;
  LAYER M3 ;
        RECT 9.32 27.955 9.6 28.325 ;
  LAYER M2 ;
        RECT 9.46 28 28.38 28.28 ;
  LAYER M3 ;
        RECT 28.24 27.955 28.52 28.325 ;
  LAYER M3 ;
        RECT 28.24 21.235 28.52 21.605 ;
  LAYER M4 ;
        RECT 28.38 21.02 30.53 21.82 ;
  LAYER M3 ;
        RECT 30.39 20.58 30.67 21.42 ;
  LAYER M2 ;
        RECT 9.3 28 9.62 28.28 ;
  LAYER M3 ;
        RECT 9.32 27.98 9.6 28.3 ;
  LAYER M2 ;
        RECT 28.22 28 28.54 28.28 ;
  LAYER M3 ;
        RECT 28.24 27.98 28.52 28.3 ;
  LAYER M2 ;
        RECT 9.3 28 9.62 28.28 ;
  LAYER M3 ;
        RECT 9.32 27.98 9.6 28.3 ;
  LAYER M2 ;
        RECT 28.22 28 28.54 28.28 ;
  LAYER M3 ;
        RECT 28.24 27.98 28.52 28.3 ;
  LAYER M2 ;
        RECT 9.3 28 9.62 28.28 ;
  LAYER M3 ;
        RECT 9.32 27.98 9.6 28.3 ;
  LAYER M2 ;
        RECT 28.22 28 28.54 28.28 ;
  LAYER M3 ;
        RECT 28.24 27.98 28.52 28.3 ;
  LAYER M3 ;
        RECT 28.24 21.235 28.52 21.605 ;
  LAYER M4 ;
        RECT 28.215 21.02 28.545 21.82 ;
  LAYER M3 ;
        RECT 30.39 21.235 30.67 21.605 ;
  LAYER M4 ;
        RECT 30.365 21.02 30.695 21.82 ;
  LAYER M2 ;
        RECT 9.3 28 9.62 28.28 ;
  LAYER M3 ;
        RECT 9.32 27.98 9.6 28.3 ;
  LAYER M2 ;
        RECT 28.22 28 28.54 28.28 ;
  LAYER M3 ;
        RECT 28.24 27.98 28.52 28.3 ;
  LAYER M3 ;
        RECT 28.24 21.235 28.52 21.605 ;
  LAYER M4 ;
        RECT 28.215 21.02 28.545 21.82 ;
  LAYER M3 ;
        RECT 30.39 21.235 30.67 21.605 ;
  LAYER M4 ;
        RECT 30.365 21.02 30.695 21.82 ;
  LAYER M3 ;
        RECT 22.22 7.82 22.5 14.02 ;
  LAYER M3 ;
        RECT 30.82 10.34 31.1 16.54 ;
  LAYER M3 ;
        RECT 31.25 2.78 31.53 7.3 ;
  LAYER M3 ;
        RECT 22.22 10.735 22.5 11.105 ;
  LAYER M2 ;
        RECT 22.36 10.78 30.96 11.06 ;
  LAYER M3 ;
        RECT 30.82 10.735 31.1 11.105 ;
  LAYER M3 ;
        RECT 30.82 7.56 31.1 10.5 ;
  LAYER M2 ;
        RECT 30.96 7.42 31.39 7.7 ;
  LAYER M3 ;
        RECT 31.25 7.14 31.53 7.56 ;
  LAYER M2 ;
        RECT 22.2 10.78 22.52 11.06 ;
  LAYER M3 ;
        RECT 22.22 10.76 22.5 11.08 ;
  LAYER M2 ;
        RECT 30.8 10.78 31.12 11.06 ;
  LAYER M3 ;
        RECT 30.82 10.76 31.1 11.08 ;
  LAYER M2 ;
        RECT 22.2 10.78 22.52 11.06 ;
  LAYER M3 ;
        RECT 22.22 10.76 22.5 11.08 ;
  LAYER M2 ;
        RECT 30.8 10.78 31.12 11.06 ;
  LAYER M3 ;
        RECT 30.82 10.76 31.1 11.08 ;
  LAYER M2 ;
        RECT 22.2 10.78 22.52 11.06 ;
  LAYER M3 ;
        RECT 22.22 10.76 22.5 11.08 ;
  LAYER M2 ;
        RECT 30.8 7.42 31.12 7.7 ;
  LAYER M3 ;
        RECT 30.82 7.4 31.1 7.72 ;
  LAYER M2 ;
        RECT 30.8 10.78 31.12 11.06 ;
  LAYER M3 ;
        RECT 30.82 10.76 31.1 11.08 ;
  LAYER M2 ;
        RECT 31.23 7.42 31.55 7.7 ;
  LAYER M3 ;
        RECT 31.25 7.4 31.53 7.72 ;
  LAYER M2 ;
        RECT 22.2 10.78 22.52 11.06 ;
  LAYER M3 ;
        RECT 22.22 10.76 22.5 11.08 ;
  LAYER M2 ;
        RECT 30.8 7.42 31.12 7.7 ;
  LAYER M3 ;
        RECT 30.82 7.4 31.1 7.72 ;
  LAYER M2 ;
        RECT 30.8 10.78 31.12 11.06 ;
  LAYER M3 ;
        RECT 30.82 10.76 31.1 11.08 ;
  LAYER M2 ;
        RECT 31.23 7.42 31.55 7.7 ;
  LAYER M3 ;
        RECT 31.25 7.4 31.53 7.72 ;
  LAYER M3 ;
        RECT 6.31 2.78 6.59 7.3 ;
  LAYER M3 ;
        RECT 6.74 10.34 7.02 16.54 ;
  LAYER M3 ;
        RECT 15.34 7.82 15.62 14.02 ;
  LAYER M3 ;
        RECT 6.31 7.14 6.59 7.56 ;
  LAYER M2 ;
        RECT 6.45 7.42 6.88 7.7 ;
  LAYER M3 ;
        RECT 6.74 7.56 7.02 10.5 ;
  LAYER M3 ;
        RECT 6.74 9.475 7.02 9.845 ;
  LAYER M2 ;
        RECT 6.88 9.52 15.48 9.8 ;
  LAYER M3 ;
        RECT 15.34 9.475 15.62 9.845 ;
  LAYER M2 ;
        RECT 6.29 7.42 6.61 7.7 ;
  LAYER M3 ;
        RECT 6.31 7.4 6.59 7.72 ;
  LAYER M2 ;
        RECT 6.72 7.42 7.04 7.7 ;
  LAYER M3 ;
        RECT 6.74 7.4 7.02 7.72 ;
  LAYER M2 ;
        RECT 6.29 7.42 6.61 7.7 ;
  LAYER M3 ;
        RECT 6.31 7.4 6.59 7.72 ;
  LAYER M2 ;
        RECT 6.72 7.42 7.04 7.7 ;
  LAYER M3 ;
        RECT 6.74 7.4 7.02 7.72 ;
  LAYER M2 ;
        RECT 6.29 7.42 6.61 7.7 ;
  LAYER M3 ;
        RECT 6.31 7.4 6.59 7.72 ;
  LAYER M2 ;
        RECT 6.72 7.42 7.04 7.7 ;
  LAYER M3 ;
        RECT 6.74 7.4 7.02 7.72 ;
  LAYER M2 ;
        RECT 6.72 9.52 7.04 9.8 ;
  LAYER M3 ;
        RECT 6.74 9.5 7.02 9.82 ;
  LAYER M2 ;
        RECT 15.32 9.52 15.64 9.8 ;
  LAYER M3 ;
        RECT 15.34 9.5 15.62 9.82 ;
  LAYER M2 ;
        RECT 6.29 7.42 6.61 7.7 ;
  LAYER M3 ;
        RECT 6.31 7.4 6.59 7.72 ;
  LAYER M2 ;
        RECT 6.72 7.42 7.04 7.7 ;
  LAYER M3 ;
        RECT 6.74 7.4 7.02 7.72 ;
  LAYER M2 ;
        RECT 6.72 9.52 7.04 9.8 ;
  LAYER M3 ;
        RECT 6.74 9.5 7.02 9.82 ;
  LAYER M2 ;
        RECT 15.32 9.52 15.64 9.8 ;
  LAYER M3 ;
        RECT 15.34 9.5 15.62 9.82 ;
  LAYER M3 ;
        RECT 16.2 8.24 16.48 14.44 ;
  LAYER M3 ;
        RECT 21.36 8.24 21.64 14.44 ;
  LAYER M2 ;
        RECT 20.04 7 28.12 7.28 ;
  LAYER M3 ;
        RECT 16.2 9.895 16.48 10.265 ;
  LAYER M2 ;
        RECT 16.34 9.94 21.5 10.22 ;
  LAYER M3 ;
        RECT 21.36 9.895 21.64 10.265 ;
  LAYER M3 ;
        RECT 21.36 7.14 21.64 8.4 ;
  LAYER M2 ;
        RECT 21.34 7 21.66 7.28 ;
  LAYER M2 ;
        RECT 16.18 9.94 16.5 10.22 ;
  LAYER M3 ;
        RECT 16.2 9.92 16.48 10.24 ;
  LAYER M2 ;
        RECT 21.34 9.94 21.66 10.22 ;
  LAYER M3 ;
        RECT 21.36 9.92 21.64 10.24 ;
  LAYER M2 ;
        RECT 16.18 9.94 16.5 10.22 ;
  LAYER M3 ;
        RECT 16.2 9.92 16.48 10.24 ;
  LAYER M2 ;
        RECT 21.34 9.94 21.66 10.22 ;
  LAYER M3 ;
        RECT 21.36 9.92 21.64 10.24 ;
  LAYER M2 ;
        RECT 16.18 9.94 16.5 10.22 ;
  LAYER M3 ;
        RECT 16.2 9.92 16.48 10.24 ;
  LAYER M2 ;
        RECT 21.34 7 21.66 7.28 ;
  LAYER M3 ;
        RECT 21.36 6.98 21.64 7.3 ;
  LAYER M2 ;
        RECT 21.34 9.94 21.66 10.22 ;
  LAYER M3 ;
        RECT 21.36 9.92 21.64 10.24 ;
  LAYER M2 ;
        RECT 16.18 9.94 16.5 10.22 ;
  LAYER M3 ;
        RECT 16.2 9.92 16.48 10.24 ;
  LAYER M2 ;
        RECT 21.34 7 21.66 7.28 ;
  LAYER M3 ;
        RECT 21.36 6.98 21.64 7.3 ;
  LAYER M2 ;
        RECT 21.34 9.94 21.66 10.22 ;
  LAYER M3 ;
        RECT 21.36 9.92 21.64 10.24 ;
  LAYER M1 ;
        RECT 17.505 3.695 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.505 2.435 17.755 3.445 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 1.345 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 9.72 2.8 17.8 3.08 ;
  LAYER M2 ;
        RECT 9.72 7 17.8 7.28 ;
  LAYER M2 ;
        RECT 9.72 0.7 17.8 0.98 ;
  LAYER M2 ;
        RECT 9.29 6.58 18.23 6.86 ;
  LAYER M3 ;
        RECT 13.62 2.78 13.9 7.3 ;
  LAYER M3 ;
        RECT 13.19 0.68 13.47 6.88 ;
  LAYER M1 ;
        RECT 36.425 21.335 36.675 24.865 ;
  LAYER M1 ;
        RECT 36.425 25.115 36.675 26.125 ;
  LAYER M1 ;
        RECT 36.425 27.215 36.675 30.745 ;
  LAYER M1 ;
        RECT 36.425 30.995 36.675 32.005 ;
  LAYER M1 ;
        RECT 36.425 33.095 36.675 36.625 ;
  LAYER M1 ;
        RECT 36.425 36.875 36.675 37.885 ;
  LAYER M1 ;
        RECT 36.425 38.975 36.675 42.505 ;
  LAYER M1 ;
        RECT 36.425 42.755 36.675 43.765 ;
  LAYER M1 ;
        RECT 36.425 44.855 36.675 45.865 ;
  LAYER M1 ;
        RECT 36.855 21.335 37.105 24.865 ;
  LAYER M1 ;
        RECT 36.855 27.215 37.105 30.745 ;
  LAYER M1 ;
        RECT 36.855 33.095 37.105 36.625 ;
  LAYER M1 ;
        RECT 36.855 38.975 37.105 42.505 ;
  LAYER M1 ;
        RECT 35.995 21.335 36.245 24.865 ;
  LAYER M1 ;
        RECT 35.995 27.215 36.245 30.745 ;
  LAYER M1 ;
        RECT 35.995 33.095 36.245 36.625 ;
  LAYER M1 ;
        RECT 35.995 38.975 36.245 42.505 ;
  LAYER M1 ;
        RECT 35.565 21.335 35.815 24.865 ;
  LAYER M1 ;
        RECT 35.565 25.115 35.815 26.125 ;
  LAYER M1 ;
        RECT 35.565 27.215 35.815 30.745 ;
  LAYER M1 ;
        RECT 35.565 30.995 35.815 32.005 ;
  LAYER M1 ;
        RECT 35.565 33.095 35.815 36.625 ;
  LAYER M1 ;
        RECT 35.565 36.875 35.815 37.885 ;
  LAYER M1 ;
        RECT 35.565 38.975 35.815 42.505 ;
  LAYER M1 ;
        RECT 35.565 42.755 35.815 43.765 ;
  LAYER M1 ;
        RECT 35.565 44.855 35.815 45.865 ;
  LAYER M1 ;
        RECT 35.135 21.335 35.385 24.865 ;
  LAYER M1 ;
        RECT 35.135 27.215 35.385 30.745 ;
  LAYER M1 ;
        RECT 35.135 33.095 35.385 36.625 ;
  LAYER M1 ;
        RECT 35.135 38.975 35.385 42.505 ;
  LAYER M1 ;
        RECT 34.705 21.335 34.955 24.865 ;
  LAYER M1 ;
        RECT 34.705 25.115 34.955 26.125 ;
  LAYER M1 ;
        RECT 34.705 27.215 34.955 30.745 ;
  LAYER M1 ;
        RECT 34.705 30.995 34.955 32.005 ;
  LAYER M1 ;
        RECT 34.705 33.095 34.955 36.625 ;
  LAYER M1 ;
        RECT 34.705 36.875 34.955 37.885 ;
  LAYER M1 ;
        RECT 34.705 38.975 34.955 42.505 ;
  LAYER M1 ;
        RECT 34.705 42.755 34.955 43.765 ;
  LAYER M1 ;
        RECT 34.705 44.855 34.955 45.865 ;
  LAYER M1 ;
        RECT 34.275 21.335 34.525 24.865 ;
  LAYER M1 ;
        RECT 34.275 27.215 34.525 30.745 ;
  LAYER M1 ;
        RECT 34.275 33.095 34.525 36.625 ;
  LAYER M1 ;
        RECT 34.275 38.975 34.525 42.505 ;
  LAYER M1 ;
        RECT 33.845 21.335 34.095 24.865 ;
  LAYER M1 ;
        RECT 33.845 25.115 34.095 26.125 ;
  LAYER M1 ;
        RECT 33.845 27.215 34.095 30.745 ;
  LAYER M1 ;
        RECT 33.845 30.995 34.095 32.005 ;
  LAYER M1 ;
        RECT 33.845 33.095 34.095 36.625 ;
  LAYER M1 ;
        RECT 33.845 36.875 34.095 37.885 ;
  LAYER M1 ;
        RECT 33.845 38.975 34.095 42.505 ;
  LAYER M1 ;
        RECT 33.845 42.755 34.095 43.765 ;
  LAYER M1 ;
        RECT 33.845 44.855 34.095 45.865 ;
  LAYER M1 ;
        RECT 33.415 21.335 33.665 24.865 ;
  LAYER M1 ;
        RECT 33.415 27.215 33.665 30.745 ;
  LAYER M1 ;
        RECT 33.415 33.095 33.665 36.625 ;
  LAYER M1 ;
        RECT 33.415 38.975 33.665 42.505 ;
  LAYER M1 ;
        RECT 32.985 21.335 33.235 24.865 ;
  LAYER M1 ;
        RECT 32.985 25.115 33.235 26.125 ;
  LAYER M1 ;
        RECT 32.985 27.215 33.235 30.745 ;
  LAYER M1 ;
        RECT 32.985 30.995 33.235 32.005 ;
  LAYER M1 ;
        RECT 32.985 33.095 33.235 36.625 ;
  LAYER M1 ;
        RECT 32.985 36.875 33.235 37.885 ;
  LAYER M1 ;
        RECT 32.985 38.975 33.235 42.505 ;
  LAYER M1 ;
        RECT 32.985 42.755 33.235 43.765 ;
  LAYER M1 ;
        RECT 32.985 44.855 33.235 45.865 ;
  LAYER M1 ;
        RECT 32.555 21.335 32.805 24.865 ;
  LAYER M1 ;
        RECT 32.555 27.215 32.805 30.745 ;
  LAYER M1 ;
        RECT 32.555 33.095 32.805 36.625 ;
  LAYER M1 ;
        RECT 32.555 38.975 32.805 42.505 ;
  LAYER M1 ;
        RECT 32.125 21.335 32.375 24.865 ;
  LAYER M1 ;
        RECT 32.125 25.115 32.375 26.125 ;
  LAYER M1 ;
        RECT 32.125 27.215 32.375 30.745 ;
  LAYER M1 ;
        RECT 32.125 30.995 32.375 32.005 ;
  LAYER M1 ;
        RECT 32.125 33.095 32.375 36.625 ;
  LAYER M1 ;
        RECT 32.125 36.875 32.375 37.885 ;
  LAYER M1 ;
        RECT 32.125 38.975 32.375 42.505 ;
  LAYER M1 ;
        RECT 32.125 42.755 32.375 43.765 ;
  LAYER M1 ;
        RECT 32.125 44.855 32.375 45.865 ;
  LAYER M1 ;
        RECT 31.695 21.335 31.945 24.865 ;
  LAYER M1 ;
        RECT 31.695 27.215 31.945 30.745 ;
  LAYER M1 ;
        RECT 31.695 33.095 31.945 36.625 ;
  LAYER M1 ;
        RECT 31.695 38.975 31.945 42.505 ;
  LAYER M1 ;
        RECT 31.265 21.335 31.515 24.865 ;
  LAYER M1 ;
        RECT 31.265 25.115 31.515 26.125 ;
  LAYER M1 ;
        RECT 31.265 27.215 31.515 30.745 ;
  LAYER M1 ;
        RECT 31.265 30.995 31.515 32.005 ;
  LAYER M1 ;
        RECT 31.265 33.095 31.515 36.625 ;
  LAYER M1 ;
        RECT 31.265 36.875 31.515 37.885 ;
  LAYER M1 ;
        RECT 31.265 38.975 31.515 42.505 ;
  LAYER M1 ;
        RECT 31.265 42.755 31.515 43.765 ;
  LAYER M1 ;
        RECT 31.265 44.855 31.515 45.865 ;
  LAYER M1 ;
        RECT 30.835 21.335 31.085 24.865 ;
  LAYER M1 ;
        RECT 30.835 27.215 31.085 30.745 ;
  LAYER M1 ;
        RECT 30.835 33.095 31.085 36.625 ;
  LAYER M1 ;
        RECT 30.835 38.975 31.085 42.505 ;
  LAYER M1 ;
        RECT 30.405 21.335 30.655 24.865 ;
  LAYER M1 ;
        RECT 30.405 25.115 30.655 26.125 ;
  LAYER M1 ;
        RECT 30.405 27.215 30.655 30.745 ;
  LAYER M1 ;
        RECT 30.405 30.995 30.655 32.005 ;
  LAYER M1 ;
        RECT 30.405 33.095 30.655 36.625 ;
  LAYER M1 ;
        RECT 30.405 36.875 30.655 37.885 ;
  LAYER M1 ;
        RECT 30.405 38.975 30.655 42.505 ;
  LAYER M1 ;
        RECT 30.405 42.755 30.655 43.765 ;
  LAYER M1 ;
        RECT 30.405 44.855 30.655 45.865 ;
  LAYER M1 ;
        RECT 29.975 21.335 30.225 24.865 ;
  LAYER M1 ;
        RECT 29.975 27.215 30.225 30.745 ;
  LAYER M1 ;
        RECT 29.975 33.095 30.225 36.625 ;
  LAYER M1 ;
        RECT 29.975 38.975 30.225 42.505 ;
  LAYER M1 ;
        RECT 29.545 21.335 29.795 24.865 ;
  LAYER M1 ;
        RECT 29.545 25.115 29.795 26.125 ;
  LAYER M1 ;
        RECT 29.545 27.215 29.795 30.745 ;
  LAYER M1 ;
        RECT 29.545 30.995 29.795 32.005 ;
  LAYER M1 ;
        RECT 29.545 33.095 29.795 36.625 ;
  LAYER M1 ;
        RECT 29.545 36.875 29.795 37.885 ;
  LAYER M1 ;
        RECT 29.545 38.975 29.795 42.505 ;
  LAYER M1 ;
        RECT 29.545 42.755 29.795 43.765 ;
  LAYER M1 ;
        RECT 29.545 44.855 29.795 45.865 ;
  LAYER M1 ;
        RECT 29.115 21.335 29.365 24.865 ;
  LAYER M1 ;
        RECT 29.115 27.215 29.365 30.745 ;
  LAYER M1 ;
        RECT 29.115 33.095 29.365 36.625 ;
  LAYER M1 ;
        RECT 29.115 38.975 29.365 42.505 ;
  LAYER M1 ;
        RECT 28.685 21.335 28.935 24.865 ;
  LAYER M1 ;
        RECT 28.685 25.115 28.935 26.125 ;
  LAYER M1 ;
        RECT 28.685 27.215 28.935 30.745 ;
  LAYER M1 ;
        RECT 28.685 30.995 28.935 32.005 ;
  LAYER M1 ;
        RECT 28.685 33.095 28.935 36.625 ;
  LAYER M1 ;
        RECT 28.685 36.875 28.935 37.885 ;
  LAYER M1 ;
        RECT 28.685 38.975 28.935 42.505 ;
  LAYER M1 ;
        RECT 28.685 42.755 28.935 43.765 ;
  LAYER M1 ;
        RECT 28.685 44.855 28.935 45.865 ;
  LAYER M1 ;
        RECT 28.255 21.335 28.505 24.865 ;
  LAYER M1 ;
        RECT 28.255 27.215 28.505 30.745 ;
  LAYER M1 ;
        RECT 28.255 33.095 28.505 36.625 ;
  LAYER M1 ;
        RECT 28.255 38.975 28.505 42.505 ;
  LAYER M1 ;
        RECT 27.825 21.335 28.075 24.865 ;
  LAYER M1 ;
        RECT 27.825 25.115 28.075 26.125 ;
  LAYER M1 ;
        RECT 27.825 27.215 28.075 30.745 ;
  LAYER M1 ;
        RECT 27.825 30.995 28.075 32.005 ;
  LAYER M1 ;
        RECT 27.825 33.095 28.075 36.625 ;
  LAYER M1 ;
        RECT 27.825 36.875 28.075 37.885 ;
  LAYER M1 ;
        RECT 27.825 38.975 28.075 42.505 ;
  LAYER M1 ;
        RECT 27.825 42.755 28.075 43.765 ;
  LAYER M1 ;
        RECT 27.825 44.855 28.075 45.865 ;
  LAYER M1 ;
        RECT 27.395 21.335 27.645 24.865 ;
  LAYER M1 ;
        RECT 27.395 27.215 27.645 30.745 ;
  LAYER M1 ;
        RECT 27.395 33.095 27.645 36.625 ;
  LAYER M1 ;
        RECT 27.395 38.975 27.645 42.505 ;
  LAYER M1 ;
        RECT 26.965 21.335 27.215 24.865 ;
  LAYER M1 ;
        RECT 26.965 25.115 27.215 26.125 ;
  LAYER M1 ;
        RECT 26.965 27.215 27.215 30.745 ;
  LAYER M1 ;
        RECT 26.965 30.995 27.215 32.005 ;
  LAYER M1 ;
        RECT 26.965 33.095 27.215 36.625 ;
  LAYER M1 ;
        RECT 26.965 36.875 27.215 37.885 ;
  LAYER M1 ;
        RECT 26.965 38.975 27.215 42.505 ;
  LAYER M1 ;
        RECT 26.965 42.755 27.215 43.765 ;
  LAYER M1 ;
        RECT 26.965 44.855 27.215 45.865 ;
  LAYER M1 ;
        RECT 26.535 21.335 26.785 24.865 ;
  LAYER M1 ;
        RECT 26.535 27.215 26.785 30.745 ;
  LAYER M1 ;
        RECT 26.535 33.095 26.785 36.625 ;
  LAYER M1 ;
        RECT 26.535 38.975 26.785 42.505 ;
  LAYER M1 ;
        RECT 26.105 21.335 26.355 24.865 ;
  LAYER M1 ;
        RECT 26.105 25.115 26.355 26.125 ;
  LAYER M1 ;
        RECT 26.105 27.215 26.355 30.745 ;
  LAYER M1 ;
        RECT 26.105 30.995 26.355 32.005 ;
  LAYER M1 ;
        RECT 26.105 33.095 26.355 36.625 ;
  LAYER M1 ;
        RECT 26.105 36.875 26.355 37.885 ;
  LAYER M1 ;
        RECT 26.105 38.975 26.355 42.505 ;
  LAYER M1 ;
        RECT 26.105 42.755 26.355 43.765 ;
  LAYER M1 ;
        RECT 26.105 44.855 26.355 45.865 ;
  LAYER M1 ;
        RECT 25.675 21.335 25.925 24.865 ;
  LAYER M1 ;
        RECT 25.675 27.215 25.925 30.745 ;
  LAYER M1 ;
        RECT 25.675 33.095 25.925 36.625 ;
  LAYER M1 ;
        RECT 25.675 38.975 25.925 42.505 ;
  LAYER M1 ;
        RECT 25.245 21.335 25.495 24.865 ;
  LAYER M1 ;
        RECT 25.245 25.115 25.495 26.125 ;
  LAYER M1 ;
        RECT 25.245 27.215 25.495 30.745 ;
  LAYER M1 ;
        RECT 25.245 30.995 25.495 32.005 ;
  LAYER M1 ;
        RECT 25.245 33.095 25.495 36.625 ;
  LAYER M1 ;
        RECT 25.245 36.875 25.495 37.885 ;
  LAYER M1 ;
        RECT 25.245 38.975 25.495 42.505 ;
  LAYER M1 ;
        RECT 25.245 42.755 25.495 43.765 ;
  LAYER M1 ;
        RECT 25.245 44.855 25.495 45.865 ;
  LAYER M1 ;
        RECT 24.815 21.335 25.065 24.865 ;
  LAYER M1 ;
        RECT 24.815 27.215 25.065 30.745 ;
  LAYER M1 ;
        RECT 24.815 33.095 25.065 36.625 ;
  LAYER M1 ;
        RECT 24.815 38.975 25.065 42.505 ;
  LAYER M1 ;
        RECT 24.385 21.335 24.635 24.865 ;
  LAYER M1 ;
        RECT 24.385 25.115 24.635 26.125 ;
  LAYER M1 ;
        RECT 24.385 27.215 24.635 30.745 ;
  LAYER M1 ;
        RECT 24.385 30.995 24.635 32.005 ;
  LAYER M1 ;
        RECT 24.385 33.095 24.635 36.625 ;
  LAYER M1 ;
        RECT 24.385 36.875 24.635 37.885 ;
  LAYER M1 ;
        RECT 24.385 38.975 24.635 42.505 ;
  LAYER M1 ;
        RECT 24.385 42.755 24.635 43.765 ;
  LAYER M1 ;
        RECT 24.385 44.855 24.635 45.865 ;
  LAYER M1 ;
        RECT 23.955 21.335 24.205 24.865 ;
  LAYER M1 ;
        RECT 23.955 27.215 24.205 30.745 ;
  LAYER M1 ;
        RECT 23.955 33.095 24.205 36.625 ;
  LAYER M1 ;
        RECT 23.955 38.975 24.205 42.505 ;
  LAYER M1 ;
        RECT 23.525 21.335 23.775 24.865 ;
  LAYER M1 ;
        RECT 23.525 25.115 23.775 26.125 ;
  LAYER M1 ;
        RECT 23.525 27.215 23.775 30.745 ;
  LAYER M1 ;
        RECT 23.525 30.995 23.775 32.005 ;
  LAYER M1 ;
        RECT 23.525 33.095 23.775 36.625 ;
  LAYER M1 ;
        RECT 23.525 36.875 23.775 37.885 ;
  LAYER M1 ;
        RECT 23.525 38.975 23.775 42.505 ;
  LAYER M1 ;
        RECT 23.525 42.755 23.775 43.765 ;
  LAYER M1 ;
        RECT 23.525 44.855 23.775 45.865 ;
  LAYER M1 ;
        RECT 23.095 21.335 23.345 24.865 ;
  LAYER M1 ;
        RECT 23.095 27.215 23.345 30.745 ;
  LAYER M1 ;
        RECT 23.095 33.095 23.345 36.625 ;
  LAYER M1 ;
        RECT 23.095 38.975 23.345 42.505 ;
  LAYER M1 ;
        RECT 22.665 21.335 22.915 24.865 ;
  LAYER M1 ;
        RECT 22.665 25.115 22.915 26.125 ;
  LAYER M1 ;
        RECT 22.665 27.215 22.915 30.745 ;
  LAYER M1 ;
        RECT 22.665 30.995 22.915 32.005 ;
  LAYER M1 ;
        RECT 22.665 33.095 22.915 36.625 ;
  LAYER M1 ;
        RECT 22.665 36.875 22.915 37.885 ;
  LAYER M1 ;
        RECT 22.665 38.975 22.915 42.505 ;
  LAYER M1 ;
        RECT 22.665 42.755 22.915 43.765 ;
  LAYER M1 ;
        RECT 22.665 44.855 22.915 45.865 ;
  LAYER M1 ;
        RECT 22.235 21.335 22.485 24.865 ;
  LAYER M1 ;
        RECT 22.235 27.215 22.485 30.745 ;
  LAYER M1 ;
        RECT 22.235 33.095 22.485 36.625 ;
  LAYER M1 ;
        RECT 22.235 38.975 22.485 42.505 ;
  LAYER M1 ;
        RECT 21.805 21.335 22.055 24.865 ;
  LAYER M1 ;
        RECT 21.805 25.115 22.055 26.125 ;
  LAYER M1 ;
        RECT 21.805 27.215 22.055 30.745 ;
  LAYER M1 ;
        RECT 21.805 30.995 22.055 32.005 ;
  LAYER M1 ;
        RECT 21.805 33.095 22.055 36.625 ;
  LAYER M1 ;
        RECT 21.805 36.875 22.055 37.885 ;
  LAYER M1 ;
        RECT 21.805 38.975 22.055 42.505 ;
  LAYER M1 ;
        RECT 21.805 42.755 22.055 43.765 ;
  LAYER M1 ;
        RECT 21.805 44.855 22.055 45.865 ;
  LAYER M1 ;
        RECT 21.375 21.335 21.625 24.865 ;
  LAYER M1 ;
        RECT 21.375 27.215 21.625 30.745 ;
  LAYER M1 ;
        RECT 21.375 33.095 21.625 36.625 ;
  LAYER M1 ;
        RECT 21.375 38.975 21.625 42.505 ;
  LAYER M1 ;
        RECT 20.945 21.335 21.195 24.865 ;
  LAYER M1 ;
        RECT 20.945 25.115 21.195 26.125 ;
  LAYER M1 ;
        RECT 20.945 27.215 21.195 30.745 ;
  LAYER M1 ;
        RECT 20.945 30.995 21.195 32.005 ;
  LAYER M1 ;
        RECT 20.945 33.095 21.195 36.625 ;
  LAYER M1 ;
        RECT 20.945 36.875 21.195 37.885 ;
  LAYER M1 ;
        RECT 20.945 38.975 21.195 42.505 ;
  LAYER M1 ;
        RECT 20.945 42.755 21.195 43.765 ;
  LAYER M1 ;
        RECT 20.945 44.855 21.195 45.865 ;
  LAYER M1 ;
        RECT 20.515 21.335 20.765 24.865 ;
  LAYER M1 ;
        RECT 20.515 27.215 20.765 30.745 ;
  LAYER M1 ;
        RECT 20.515 33.095 20.765 36.625 ;
  LAYER M1 ;
        RECT 20.515 38.975 20.765 42.505 ;
  LAYER M1 ;
        RECT 20.085 21.335 20.335 24.865 ;
  LAYER M1 ;
        RECT 20.085 25.115 20.335 26.125 ;
  LAYER M1 ;
        RECT 20.085 27.215 20.335 30.745 ;
  LAYER M1 ;
        RECT 20.085 30.995 20.335 32.005 ;
  LAYER M1 ;
        RECT 20.085 33.095 20.335 36.625 ;
  LAYER M1 ;
        RECT 20.085 36.875 20.335 37.885 ;
  LAYER M1 ;
        RECT 20.085 38.975 20.335 42.505 ;
  LAYER M1 ;
        RECT 20.085 42.755 20.335 43.765 ;
  LAYER M1 ;
        RECT 20.085 44.855 20.335 45.865 ;
  LAYER M1 ;
        RECT 19.655 21.335 19.905 24.865 ;
  LAYER M1 ;
        RECT 19.655 27.215 19.905 30.745 ;
  LAYER M1 ;
        RECT 19.655 33.095 19.905 36.625 ;
  LAYER M1 ;
        RECT 19.655 38.975 19.905 42.505 ;
  LAYER M2 ;
        RECT 20.04 25.48 36.72 25.76 ;
  LAYER M2 ;
        RECT 20.04 21.28 36.72 21.56 ;
  LAYER M2 ;
        RECT 19.61 21.7 37.15 21.98 ;
  LAYER M2 ;
        RECT 20.04 31.36 36.72 31.64 ;
  LAYER M2 ;
        RECT 20.04 27.16 36.72 27.44 ;
  LAYER M2 ;
        RECT 19.61 27.58 37.15 27.86 ;
  LAYER M2 ;
        RECT 20.04 37.24 36.72 37.52 ;
  LAYER M2 ;
        RECT 20.04 33.04 36.72 33.32 ;
  LAYER M2 ;
        RECT 19.61 33.46 37.15 33.74 ;
  LAYER M2 ;
        RECT 20.04 43.12 36.72 43.4 ;
  LAYER M2 ;
        RECT 20.04 38.92 36.72 39.2 ;
  LAYER M2 ;
        RECT 20.04 45.22 36.72 45.5 ;
  LAYER M2 ;
        RECT 19.61 39.34 37.15 39.62 ;
  LAYER M3 ;
        RECT 28.24 21.26 28.52 43.42 ;
  LAYER M3 ;
        RECT 27.81 21.68 28.09 45.52 ;
  LAYER M1 ;
        RECT 32.125 3.695 32.375 7.225 ;
  LAYER M1 ;
        RECT 32.125 2.435 32.375 3.445 ;
  LAYER M1 ;
        RECT 32.125 0.335 32.375 1.345 ;
  LAYER M1 ;
        RECT 32.555 3.695 32.805 7.225 ;
  LAYER M1 ;
        RECT 31.695 3.695 31.945 7.225 ;
  LAYER M1 ;
        RECT 31.265 3.695 31.515 7.225 ;
  LAYER M1 ;
        RECT 31.265 2.435 31.515 3.445 ;
  LAYER M1 ;
        RECT 31.265 0.335 31.515 1.345 ;
  LAYER M1 ;
        RECT 30.835 3.695 31.085 7.225 ;
  LAYER M1 ;
        RECT 30.405 3.695 30.655 7.225 ;
  LAYER M1 ;
        RECT 30.405 2.435 30.655 3.445 ;
  LAYER M1 ;
        RECT 30.405 0.335 30.655 1.345 ;
  LAYER M1 ;
        RECT 29.975 3.695 30.225 7.225 ;
  LAYER M2 ;
        RECT 30.36 2.8 32.42 3.08 ;
  LAYER M2 ;
        RECT 30.36 7 32.42 7.28 ;
  LAYER M2 ;
        RECT 30.36 0.7 32.42 0.98 ;
  LAYER M2 ;
        RECT 29.93 6.58 32.85 6.86 ;
  LAYER M3 ;
        RECT 31.25 2.78 31.53 7.3 ;
  LAYER M3 ;
        RECT 30.82 0.68 31.1 6.88 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M2 ;
        RECT 5.42 2.8 7.48 3.08 ;
  LAYER M2 ;
        RECT 5.42 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 5.42 0.7 7.48 0.98 ;
  LAYER M2 ;
        RECT 4.99 6.58 7.91 6.86 ;
  LAYER M3 ;
        RECT 6.31 2.78 6.59 7.3 ;
  LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
  LAYER M1 ;
        RECT 1.165 21.335 1.415 24.865 ;
  LAYER M1 ;
        RECT 1.165 25.115 1.415 26.125 ;
  LAYER M1 ;
        RECT 1.165 27.215 1.415 30.745 ;
  LAYER M1 ;
        RECT 1.165 30.995 1.415 32.005 ;
  LAYER M1 ;
        RECT 1.165 33.095 1.415 36.625 ;
  LAYER M1 ;
        RECT 1.165 36.875 1.415 37.885 ;
  LAYER M1 ;
        RECT 1.165 38.975 1.415 42.505 ;
  LAYER M1 ;
        RECT 1.165 42.755 1.415 43.765 ;
  LAYER M1 ;
        RECT 1.165 44.855 1.415 45.865 ;
  LAYER M1 ;
        RECT 0.735 21.335 0.985 24.865 ;
  LAYER M1 ;
        RECT 0.735 27.215 0.985 30.745 ;
  LAYER M1 ;
        RECT 0.735 33.095 0.985 36.625 ;
  LAYER M1 ;
        RECT 0.735 38.975 0.985 42.505 ;
  LAYER M1 ;
        RECT 1.595 21.335 1.845 24.865 ;
  LAYER M1 ;
        RECT 1.595 27.215 1.845 30.745 ;
  LAYER M1 ;
        RECT 1.595 33.095 1.845 36.625 ;
  LAYER M1 ;
        RECT 1.595 38.975 1.845 42.505 ;
  LAYER M1 ;
        RECT 2.025 21.335 2.275 24.865 ;
  LAYER M1 ;
        RECT 2.025 25.115 2.275 26.125 ;
  LAYER M1 ;
        RECT 2.025 27.215 2.275 30.745 ;
  LAYER M1 ;
        RECT 2.025 30.995 2.275 32.005 ;
  LAYER M1 ;
        RECT 2.025 33.095 2.275 36.625 ;
  LAYER M1 ;
        RECT 2.025 36.875 2.275 37.885 ;
  LAYER M1 ;
        RECT 2.025 38.975 2.275 42.505 ;
  LAYER M1 ;
        RECT 2.025 42.755 2.275 43.765 ;
  LAYER M1 ;
        RECT 2.025 44.855 2.275 45.865 ;
  LAYER M1 ;
        RECT 2.455 21.335 2.705 24.865 ;
  LAYER M1 ;
        RECT 2.455 27.215 2.705 30.745 ;
  LAYER M1 ;
        RECT 2.455 33.095 2.705 36.625 ;
  LAYER M1 ;
        RECT 2.455 38.975 2.705 42.505 ;
  LAYER M1 ;
        RECT 2.885 21.335 3.135 24.865 ;
  LAYER M1 ;
        RECT 2.885 25.115 3.135 26.125 ;
  LAYER M1 ;
        RECT 2.885 27.215 3.135 30.745 ;
  LAYER M1 ;
        RECT 2.885 30.995 3.135 32.005 ;
  LAYER M1 ;
        RECT 2.885 33.095 3.135 36.625 ;
  LAYER M1 ;
        RECT 2.885 36.875 3.135 37.885 ;
  LAYER M1 ;
        RECT 2.885 38.975 3.135 42.505 ;
  LAYER M1 ;
        RECT 2.885 42.755 3.135 43.765 ;
  LAYER M1 ;
        RECT 2.885 44.855 3.135 45.865 ;
  LAYER M1 ;
        RECT 3.315 21.335 3.565 24.865 ;
  LAYER M1 ;
        RECT 3.315 27.215 3.565 30.745 ;
  LAYER M1 ;
        RECT 3.315 33.095 3.565 36.625 ;
  LAYER M1 ;
        RECT 3.315 38.975 3.565 42.505 ;
  LAYER M1 ;
        RECT 3.745 21.335 3.995 24.865 ;
  LAYER M1 ;
        RECT 3.745 25.115 3.995 26.125 ;
  LAYER M1 ;
        RECT 3.745 27.215 3.995 30.745 ;
  LAYER M1 ;
        RECT 3.745 30.995 3.995 32.005 ;
  LAYER M1 ;
        RECT 3.745 33.095 3.995 36.625 ;
  LAYER M1 ;
        RECT 3.745 36.875 3.995 37.885 ;
  LAYER M1 ;
        RECT 3.745 38.975 3.995 42.505 ;
  LAYER M1 ;
        RECT 3.745 42.755 3.995 43.765 ;
  LAYER M1 ;
        RECT 3.745 44.855 3.995 45.865 ;
  LAYER M1 ;
        RECT 4.175 21.335 4.425 24.865 ;
  LAYER M1 ;
        RECT 4.175 27.215 4.425 30.745 ;
  LAYER M1 ;
        RECT 4.175 33.095 4.425 36.625 ;
  LAYER M1 ;
        RECT 4.175 38.975 4.425 42.505 ;
  LAYER M1 ;
        RECT 4.605 21.335 4.855 24.865 ;
  LAYER M1 ;
        RECT 4.605 25.115 4.855 26.125 ;
  LAYER M1 ;
        RECT 4.605 27.215 4.855 30.745 ;
  LAYER M1 ;
        RECT 4.605 30.995 4.855 32.005 ;
  LAYER M1 ;
        RECT 4.605 33.095 4.855 36.625 ;
  LAYER M1 ;
        RECT 4.605 36.875 4.855 37.885 ;
  LAYER M1 ;
        RECT 4.605 38.975 4.855 42.505 ;
  LAYER M1 ;
        RECT 4.605 42.755 4.855 43.765 ;
  LAYER M1 ;
        RECT 4.605 44.855 4.855 45.865 ;
  LAYER M1 ;
        RECT 5.035 21.335 5.285 24.865 ;
  LAYER M1 ;
        RECT 5.035 27.215 5.285 30.745 ;
  LAYER M1 ;
        RECT 5.035 33.095 5.285 36.625 ;
  LAYER M1 ;
        RECT 5.035 38.975 5.285 42.505 ;
  LAYER M1 ;
        RECT 5.465 21.335 5.715 24.865 ;
  LAYER M1 ;
        RECT 5.465 25.115 5.715 26.125 ;
  LAYER M1 ;
        RECT 5.465 27.215 5.715 30.745 ;
  LAYER M1 ;
        RECT 5.465 30.995 5.715 32.005 ;
  LAYER M1 ;
        RECT 5.465 33.095 5.715 36.625 ;
  LAYER M1 ;
        RECT 5.465 36.875 5.715 37.885 ;
  LAYER M1 ;
        RECT 5.465 38.975 5.715 42.505 ;
  LAYER M1 ;
        RECT 5.465 42.755 5.715 43.765 ;
  LAYER M1 ;
        RECT 5.465 44.855 5.715 45.865 ;
  LAYER M1 ;
        RECT 5.895 21.335 6.145 24.865 ;
  LAYER M1 ;
        RECT 5.895 27.215 6.145 30.745 ;
  LAYER M1 ;
        RECT 5.895 33.095 6.145 36.625 ;
  LAYER M1 ;
        RECT 5.895 38.975 6.145 42.505 ;
  LAYER M1 ;
        RECT 6.325 21.335 6.575 24.865 ;
  LAYER M1 ;
        RECT 6.325 25.115 6.575 26.125 ;
  LAYER M1 ;
        RECT 6.325 27.215 6.575 30.745 ;
  LAYER M1 ;
        RECT 6.325 30.995 6.575 32.005 ;
  LAYER M1 ;
        RECT 6.325 33.095 6.575 36.625 ;
  LAYER M1 ;
        RECT 6.325 36.875 6.575 37.885 ;
  LAYER M1 ;
        RECT 6.325 38.975 6.575 42.505 ;
  LAYER M1 ;
        RECT 6.325 42.755 6.575 43.765 ;
  LAYER M1 ;
        RECT 6.325 44.855 6.575 45.865 ;
  LAYER M1 ;
        RECT 6.755 21.335 7.005 24.865 ;
  LAYER M1 ;
        RECT 6.755 27.215 7.005 30.745 ;
  LAYER M1 ;
        RECT 6.755 33.095 7.005 36.625 ;
  LAYER M1 ;
        RECT 6.755 38.975 7.005 42.505 ;
  LAYER M1 ;
        RECT 7.185 21.335 7.435 24.865 ;
  LAYER M1 ;
        RECT 7.185 25.115 7.435 26.125 ;
  LAYER M1 ;
        RECT 7.185 27.215 7.435 30.745 ;
  LAYER M1 ;
        RECT 7.185 30.995 7.435 32.005 ;
  LAYER M1 ;
        RECT 7.185 33.095 7.435 36.625 ;
  LAYER M1 ;
        RECT 7.185 36.875 7.435 37.885 ;
  LAYER M1 ;
        RECT 7.185 38.975 7.435 42.505 ;
  LAYER M1 ;
        RECT 7.185 42.755 7.435 43.765 ;
  LAYER M1 ;
        RECT 7.185 44.855 7.435 45.865 ;
  LAYER M1 ;
        RECT 7.615 21.335 7.865 24.865 ;
  LAYER M1 ;
        RECT 7.615 27.215 7.865 30.745 ;
  LAYER M1 ;
        RECT 7.615 33.095 7.865 36.625 ;
  LAYER M1 ;
        RECT 7.615 38.975 7.865 42.505 ;
  LAYER M1 ;
        RECT 8.045 21.335 8.295 24.865 ;
  LAYER M1 ;
        RECT 8.045 25.115 8.295 26.125 ;
  LAYER M1 ;
        RECT 8.045 27.215 8.295 30.745 ;
  LAYER M1 ;
        RECT 8.045 30.995 8.295 32.005 ;
  LAYER M1 ;
        RECT 8.045 33.095 8.295 36.625 ;
  LAYER M1 ;
        RECT 8.045 36.875 8.295 37.885 ;
  LAYER M1 ;
        RECT 8.045 38.975 8.295 42.505 ;
  LAYER M1 ;
        RECT 8.045 42.755 8.295 43.765 ;
  LAYER M1 ;
        RECT 8.045 44.855 8.295 45.865 ;
  LAYER M1 ;
        RECT 8.475 21.335 8.725 24.865 ;
  LAYER M1 ;
        RECT 8.475 27.215 8.725 30.745 ;
  LAYER M1 ;
        RECT 8.475 33.095 8.725 36.625 ;
  LAYER M1 ;
        RECT 8.475 38.975 8.725 42.505 ;
  LAYER M1 ;
        RECT 8.905 21.335 9.155 24.865 ;
  LAYER M1 ;
        RECT 8.905 25.115 9.155 26.125 ;
  LAYER M1 ;
        RECT 8.905 27.215 9.155 30.745 ;
  LAYER M1 ;
        RECT 8.905 30.995 9.155 32.005 ;
  LAYER M1 ;
        RECT 8.905 33.095 9.155 36.625 ;
  LAYER M1 ;
        RECT 8.905 36.875 9.155 37.885 ;
  LAYER M1 ;
        RECT 8.905 38.975 9.155 42.505 ;
  LAYER M1 ;
        RECT 8.905 42.755 9.155 43.765 ;
  LAYER M1 ;
        RECT 8.905 44.855 9.155 45.865 ;
  LAYER M1 ;
        RECT 9.335 21.335 9.585 24.865 ;
  LAYER M1 ;
        RECT 9.335 27.215 9.585 30.745 ;
  LAYER M1 ;
        RECT 9.335 33.095 9.585 36.625 ;
  LAYER M1 ;
        RECT 9.335 38.975 9.585 42.505 ;
  LAYER M1 ;
        RECT 9.765 21.335 10.015 24.865 ;
  LAYER M1 ;
        RECT 9.765 25.115 10.015 26.125 ;
  LAYER M1 ;
        RECT 9.765 27.215 10.015 30.745 ;
  LAYER M1 ;
        RECT 9.765 30.995 10.015 32.005 ;
  LAYER M1 ;
        RECT 9.765 33.095 10.015 36.625 ;
  LAYER M1 ;
        RECT 9.765 36.875 10.015 37.885 ;
  LAYER M1 ;
        RECT 9.765 38.975 10.015 42.505 ;
  LAYER M1 ;
        RECT 9.765 42.755 10.015 43.765 ;
  LAYER M1 ;
        RECT 9.765 44.855 10.015 45.865 ;
  LAYER M1 ;
        RECT 10.195 21.335 10.445 24.865 ;
  LAYER M1 ;
        RECT 10.195 27.215 10.445 30.745 ;
  LAYER M1 ;
        RECT 10.195 33.095 10.445 36.625 ;
  LAYER M1 ;
        RECT 10.195 38.975 10.445 42.505 ;
  LAYER M1 ;
        RECT 10.625 21.335 10.875 24.865 ;
  LAYER M1 ;
        RECT 10.625 25.115 10.875 26.125 ;
  LAYER M1 ;
        RECT 10.625 27.215 10.875 30.745 ;
  LAYER M1 ;
        RECT 10.625 30.995 10.875 32.005 ;
  LAYER M1 ;
        RECT 10.625 33.095 10.875 36.625 ;
  LAYER M1 ;
        RECT 10.625 36.875 10.875 37.885 ;
  LAYER M1 ;
        RECT 10.625 38.975 10.875 42.505 ;
  LAYER M1 ;
        RECT 10.625 42.755 10.875 43.765 ;
  LAYER M1 ;
        RECT 10.625 44.855 10.875 45.865 ;
  LAYER M1 ;
        RECT 11.055 21.335 11.305 24.865 ;
  LAYER M1 ;
        RECT 11.055 27.215 11.305 30.745 ;
  LAYER M1 ;
        RECT 11.055 33.095 11.305 36.625 ;
  LAYER M1 ;
        RECT 11.055 38.975 11.305 42.505 ;
  LAYER M1 ;
        RECT 11.485 21.335 11.735 24.865 ;
  LAYER M1 ;
        RECT 11.485 25.115 11.735 26.125 ;
  LAYER M1 ;
        RECT 11.485 27.215 11.735 30.745 ;
  LAYER M1 ;
        RECT 11.485 30.995 11.735 32.005 ;
  LAYER M1 ;
        RECT 11.485 33.095 11.735 36.625 ;
  LAYER M1 ;
        RECT 11.485 36.875 11.735 37.885 ;
  LAYER M1 ;
        RECT 11.485 38.975 11.735 42.505 ;
  LAYER M1 ;
        RECT 11.485 42.755 11.735 43.765 ;
  LAYER M1 ;
        RECT 11.485 44.855 11.735 45.865 ;
  LAYER M1 ;
        RECT 11.915 21.335 12.165 24.865 ;
  LAYER M1 ;
        RECT 11.915 27.215 12.165 30.745 ;
  LAYER M1 ;
        RECT 11.915 33.095 12.165 36.625 ;
  LAYER M1 ;
        RECT 11.915 38.975 12.165 42.505 ;
  LAYER M1 ;
        RECT 12.345 21.335 12.595 24.865 ;
  LAYER M1 ;
        RECT 12.345 25.115 12.595 26.125 ;
  LAYER M1 ;
        RECT 12.345 27.215 12.595 30.745 ;
  LAYER M1 ;
        RECT 12.345 30.995 12.595 32.005 ;
  LAYER M1 ;
        RECT 12.345 33.095 12.595 36.625 ;
  LAYER M1 ;
        RECT 12.345 36.875 12.595 37.885 ;
  LAYER M1 ;
        RECT 12.345 38.975 12.595 42.505 ;
  LAYER M1 ;
        RECT 12.345 42.755 12.595 43.765 ;
  LAYER M1 ;
        RECT 12.345 44.855 12.595 45.865 ;
  LAYER M1 ;
        RECT 12.775 21.335 13.025 24.865 ;
  LAYER M1 ;
        RECT 12.775 27.215 13.025 30.745 ;
  LAYER M1 ;
        RECT 12.775 33.095 13.025 36.625 ;
  LAYER M1 ;
        RECT 12.775 38.975 13.025 42.505 ;
  LAYER M1 ;
        RECT 13.205 21.335 13.455 24.865 ;
  LAYER M1 ;
        RECT 13.205 25.115 13.455 26.125 ;
  LAYER M1 ;
        RECT 13.205 27.215 13.455 30.745 ;
  LAYER M1 ;
        RECT 13.205 30.995 13.455 32.005 ;
  LAYER M1 ;
        RECT 13.205 33.095 13.455 36.625 ;
  LAYER M1 ;
        RECT 13.205 36.875 13.455 37.885 ;
  LAYER M1 ;
        RECT 13.205 38.975 13.455 42.505 ;
  LAYER M1 ;
        RECT 13.205 42.755 13.455 43.765 ;
  LAYER M1 ;
        RECT 13.205 44.855 13.455 45.865 ;
  LAYER M1 ;
        RECT 13.635 21.335 13.885 24.865 ;
  LAYER M1 ;
        RECT 13.635 27.215 13.885 30.745 ;
  LAYER M1 ;
        RECT 13.635 33.095 13.885 36.625 ;
  LAYER M1 ;
        RECT 13.635 38.975 13.885 42.505 ;
  LAYER M1 ;
        RECT 14.065 21.335 14.315 24.865 ;
  LAYER M1 ;
        RECT 14.065 25.115 14.315 26.125 ;
  LAYER M1 ;
        RECT 14.065 27.215 14.315 30.745 ;
  LAYER M1 ;
        RECT 14.065 30.995 14.315 32.005 ;
  LAYER M1 ;
        RECT 14.065 33.095 14.315 36.625 ;
  LAYER M1 ;
        RECT 14.065 36.875 14.315 37.885 ;
  LAYER M1 ;
        RECT 14.065 38.975 14.315 42.505 ;
  LAYER M1 ;
        RECT 14.065 42.755 14.315 43.765 ;
  LAYER M1 ;
        RECT 14.065 44.855 14.315 45.865 ;
  LAYER M1 ;
        RECT 14.495 21.335 14.745 24.865 ;
  LAYER M1 ;
        RECT 14.495 27.215 14.745 30.745 ;
  LAYER M1 ;
        RECT 14.495 33.095 14.745 36.625 ;
  LAYER M1 ;
        RECT 14.495 38.975 14.745 42.505 ;
  LAYER M1 ;
        RECT 14.925 21.335 15.175 24.865 ;
  LAYER M1 ;
        RECT 14.925 25.115 15.175 26.125 ;
  LAYER M1 ;
        RECT 14.925 27.215 15.175 30.745 ;
  LAYER M1 ;
        RECT 14.925 30.995 15.175 32.005 ;
  LAYER M1 ;
        RECT 14.925 33.095 15.175 36.625 ;
  LAYER M1 ;
        RECT 14.925 36.875 15.175 37.885 ;
  LAYER M1 ;
        RECT 14.925 38.975 15.175 42.505 ;
  LAYER M1 ;
        RECT 14.925 42.755 15.175 43.765 ;
  LAYER M1 ;
        RECT 14.925 44.855 15.175 45.865 ;
  LAYER M1 ;
        RECT 15.355 21.335 15.605 24.865 ;
  LAYER M1 ;
        RECT 15.355 27.215 15.605 30.745 ;
  LAYER M1 ;
        RECT 15.355 33.095 15.605 36.625 ;
  LAYER M1 ;
        RECT 15.355 38.975 15.605 42.505 ;
  LAYER M1 ;
        RECT 15.785 21.335 16.035 24.865 ;
  LAYER M1 ;
        RECT 15.785 25.115 16.035 26.125 ;
  LAYER M1 ;
        RECT 15.785 27.215 16.035 30.745 ;
  LAYER M1 ;
        RECT 15.785 30.995 16.035 32.005 ;
  LAYER M1 ;
        RECT 15.785 33.095 16.035 36.625 ;
  LAYER M1 ;
        RECT 15.785 36.875 16.035 37.885 ;
  LAYER M1 ;
        RECT 15.785 38.975 16.035 42.505 ;
  LAYER M1 ;
        RECT 15.785 42.755 16.035 43.765 ;
  LAYER M1 ;
        RECT 15.785 44.855 16.035 45.865 ;
  LAYER M1 ;
        RECT 16.215 21.335 16.465 24.865 ;
  LAYER M1 ;
        RECT 16.215 27.215 16.465 30.745 ;
  LAYER M1 ;
        RECT 16.215 33.095 16.465 36.625 ;
  LAYER M1 ;
        RECT 16.215 38.975 16.465 42.505 ;
  LAYER M1 ;
        RECT 16.645 21.335 16.895 24.865 ;
  LAYER M1 ;
        RECT 16.645 25.115 16.895 26.125 ;
  LAYER M1 ;
        RECT 16.645 27.215 16.895 30.745 ;
  LAYER M1 ;
        RECT 16.645 30.995 16.895 32.005 ;
  LAYER M1 ;
        RECT 16.645 33.095 16.895 36.625 ;
  LAYER M1 ;
        RECT 16.645 36.875 16.895 37.885 ;
  LAYER M1 ;
        RECT 16.645 38.975 16.895 42.505 ;
  LAYER M1 ;
        RECT 16.645 42.755 16.895 43.765 ;
  LAYER M1 ;
        RECT 16.645 44.855 16.895 45.865 ;
  LAYER M1 ;
        RECT 17.075 21.335 17.325 24.865 ;
  LAYER M1 ;
        RECT 17.075 27.215 17.325 30.745 ;
  LAYER M1 ;
        RECT 17.075 33.095 17.325 36.625 ;
  LAYER M1 ;
        RECT 17.075 38.975 17.325 42.505 ;
  LAYER M1 ;
        RECT 17.505 21.335 17.755 24.865 ;
  LAYER M1 ;
        RECT 17.505 25.115 17.755 26.125 ;
  LAYER M1 ;
        RECT 17.505 27.215 17.755 30.745 ;
  LAYER M1 ;
        RECT 17.505 30.995 17.755 32.005 ;
  LAYER M1 ;
        RECT 17.505 33.095 17.755 36.625 ;
  LAYER M1 ;
        RECT 17.505 36.875 17.755 37.885 ;
  LAYER M1 ;
        RECT 17.505 38.975 17.755 42.505 ;
  LAYER M1 ;
        RECT 17.505 42.755 17.755 43.765 ;
  LAYER M1 ;
        RECT 17.505 44.855 17.755 45.865 ;
  LAYER M1 ;
        RECT 17.935 21.335 18.185 24.865 ;
  LAYER M1 ;
        RECT 17.935 27.215 18.185 30.745 ;
  LAYER M1 ;
        RECT 17.935 33.095 18.185 36.625 ;
  LAYER M1 ;
        RECT 17.935 38.975 18.185 42.505 ;
  LAYER M2 ;
        RECT 1.12 21.28 17.8 21.56 ;
  LAYER M2 ;
        RECT 1.12 25.48 17.8 25.76 ;
  LAYER M2 ;
        RECT 0.69 21.7 18.23 21.98 ;
  LAYER M2 ;
        RECT 1.12 27.16 17.8 27.44 ;
  LAYER M2 ;
        RECT 1.12 31.36 17.8 31.64 ;
  LAYER M2 ;
        RECT 0.69 27.58 18.23 27.86 ;
  LAYER M2 ;
        RECT 1.12 33.04 17.8 33.32 ;
  LAYER M2 ;
        RECT 1.12 37.24 17.8 37.52 ;
  LAYER M2 ;
        RECT 0.69 33.46 18.23 33.74 ;
  LAYER M2 ;
        RECT 1.12 38.92 17.8 39.2 ;
  LAYER M2 ;
        RECT 1.12 43.12 17.8 43.4 ;
  LAYER M2 ;
        RECT 1.12 45.22 17.8 45.5 ;
  LAYER M2 ;
        RECT 0.69 39.34 18.23 39.62 ;
  LAYER M3 ;
        RECT 8.89 21.26 9.17 39.22 ;
  LAYER M3 ;
        RECT 9.32 25.46 9.6 43.42 ;
  LAYER M3 ;
        RECT 9.75 21.68 10.03 45.52 ;
  LAYER M1 ;
        RECT 20.085 3.695 20.335 7.225 ;
  LAYER M1 ;
        RECT 20.085 2.435 20.335 3.445 ;
  LAYER M1 ;
        RECT 20.085 0.335 20.335 1.345 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M1 ;
        RECT 20.515 3.695 20.765 7.225 ;
  LAYER M1 ;
        RECT 20.945 3.695 21.195 7.225 ;
  LAYER M1 ;
        RECT 20.945 2.435 21.195 3.445 ;
  LAYER M1 ;
        RECT 20.945 0.335 21.195 1.345 ;
  LAYER M1 ;
        RECT 21.375 3.695 21.625 7.225 ;
  LAYER M1 ;
        RECT 21.805 3.695 22.055 7.225 ;
  LAYER M1 ;
        RECT 21.805 2.435 22.055 3.445 ;
  LAYER M1 ;
        RECT 21.805 0.335 22.055 1.345 ;
  LAYER M1 ;
        RECT 22.235 3.695 22.485 7.225 ;
  LAYER M1 ;
        RECT 22.665 3.695 22.915 7.225 ;
  LAYER M1 ;
        RECT 22.665 2.435 22.915 3.445 ;
  LAYER M1 ;
        RECT 22.665 0.335 22.915 1.345 ;
  LAYER M1 ;
        RECT 23.095 3.695 23.345 7.225 ;
  LAYER M1 ;
        RECT 23.525 3.695 23.775 7.225 ;
  LAYER M1 ;
        RECT 23.525 2.435 23.775 3.445 ;
  LAYER M1 ;
        RECT 23.525 0.335 23.775 1.345 ;
  LAYER M1 ;
        RECT 23.955 3.695 24.205 7.225 ;
  LAYER M1 ;
        RECT 24.385 3.695 24.635 7.225 ;
  LAYER M1 ;
        RECT 24.385 2.435 24.635 3.445 ;
  LAYER M1 ;
        RECT 24.385 0.335 24.635 1.345 ;
  LAYER M1 ;
        RECT 24.815 3.695 25.065 7.225 ;
  LAYER M1 ;
        RECT 25.245 3.695 25.495 7.225 ;
  LAYER M1 ;
        RECT 25.245 2.435 25.495 3.445 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 1.345 ;
  LAYER M1 ;
        RECT 25.675 3.695 25.925 7.225 ;
  LAYER M1 ;
        RECT 26.105 3.695 26.355 7.225 ;
  LAYER M1 ;
        RECT 26.105 2.435 26.355 3.445 ;
  LAYER M1 ;
        RECT 26.105 0.335 26.355 1.345 ;
  LAYER M1 ;
        RECT 26.535 3.695 26.785 7.225 ;
  LAYER M1 ;
        RECT 26.965 3.695 27.215 7.225 ;
  LAYER M1 ;
        RECT 26.965 2.435 27.215 3.445 ;
  LAYER M1 ;
        RECT 26.965 0.335 27.215 1.345 ;
  LAYER M1 ;
        RECT 27.395 3.695 27.645 7.225 ;
  LAYER M1 ;
        RECT 27.825 3.695 28.075 7.225 ;
  LAYER M1 ;
        RECT 27.825 2.435 28.075 3.445 ;
  LAYER M1 ;
        RECT 27.825 0.335 28.075 1.345 ;
  LAYER M1 ;
        RECT 28.255 3.695 28.505 7.225 ;
  LAYER M2 ;
        RECT 20.04 0.7 28.12 0.98 ;
  LAYER M2 ;
        RECT 19.61 6.58 28.55 6.86 ;
  LAYER M2 ;
        RECT 20.04 7 28.12 7.28 ;
  LAYER M2 ;
        RECT 20.04 2.8 28.12 3.08 ;
  LAYER M3 ;
        RECT 24.37 0.68 24.65 6.88 ;
  LAYER M1 ;
        RECT 26.105 17.135 26.355 20.665 ;
  LAYER M1 ;
        RECT 26.105 15.875 26.355 16.885 ;
  LAYER M1 ;
        RECT 26.105 11.255 26.355 14.785 ;
  LAYER M1 ;
        RECT 26.105 9.995 26.355 11.005 ;
  LAYER M1 ;
        RECT 26.105 7.895 26.355 8.905 ;
  LAYER M1 ;
        RECT 25.675 17.135 25.925 20.665 ;
  LAYER M1 ;
        RECT 25.675 11.255 25.925 14.785 ;
  LAYER M1 ;
        RECT 26.535 17.135 26.785 20.665 ;
  LAYER M1 ;
        RECT 26.535 11.255 26.785 14.785 ;
  LAYER M1 ;
        RECT 26.965 17.135 27.215 20.665 ;
  LAYER M1 ;
        RECT 26.965 15.875 27.215 16.885 ;
  LAYER M1 ;
        RECT 26.965 11.255 27.215 14.785 ;
  LAYER M1 ;
        RECT 26.965 9.995 27.215 11.005 ;
  LAYER M1 ;
        RECT 26.965 7.895 27.215 8.905 ;
  LAYER M1 ;
        RECT 27.395 17.135 27.645 20.665 ;
  LAYER M1 ;
        RECT 27.395 11.255 27.645 14.785 ;
  LAYER M1 ;
        RECT 27.825 17.135 28.075 20.665 ;
  LAYER M1 ;
        RECT 27.825 15.875 28.075 16.885 ;
  LAYER M1 ;
        RECT 27.825 11.255 28.075 14.785 ;
  LAYER M1 ;
        RECT 27.825 9.995 28.075 11.005 ;
  LAYER M1 ;
        RECT 27.825 7.895 28.075 8.905 ;
  LAYER M1 ;
        RECT 28.255 17.135 28.505 20.665 ;
  LAYER M1 ;
        RECT 28.255 11.255 28.505 14.785 ;
  LAYER M1 ;
        RECT 28.685 17.135 28.935 20.665 ;
  LAYER M1 ;
        RECT 28.685 15.875 28.935 16.885 ;
  LAYER M1 ;
        RECT 28.685 11.255 28.935 14.785 ;
  LAYER M1 ;
        RECT 28.685 9.995 28.935 11.005 ;
  LAYER M1 ;
        RECT 28.685 7.895 28.935 8.905 ;
  LAYER M1 ;
        RECT 29.115 17.135 29.365 20.665 ;
  LAYER M1 ;
        RECT 29.115 11.255 29.365 14.785 ;
  LAYER M1 ;
        RECT 29.545 17.135 29.795 20.665 ;
  LAYER M1 ;
        RECT 29.545 15.875 29.795 16.885 ;
  LAYER M1 ;
        RECT 29.545 11.255 29.795 14.785 ;
  LAYER M1 ;
        RECT 29.545 9.995 29.795 11.005 ;
  LAYER M1 ;
        RECT 29.545 7.895 29.795 8.905 ;
  LAYER M1 ;
        RECT 29.975 17.135 30.225 20.665 ;
  LAYER M1 ;
        RECT 29.975 11.255 30.225 14.785 ;
  LAYER M1 ;
        RECT 30.405 17.135 30.655 20.665 ;
  LAYER M1 ;
        RECT 30.405 15.875 30.655 16.885 ;
  LAYER M1 ;
        RECT 30.405 11.255 30.655 14.785 ;
  LAYER M1 ;
        RECT 30.405 9.995 30.655 11.005 ;
  LAYER M1 ;
        RECT 30.405 7.895 30.655 8.905 ;
  LAYER M1 ;
        RECT 30.835 17.135 31.085 20.665 ;
  LAYER M1 ;
        RECT 30.835 11.255 31.085 14.785 ;
  LAYER M1 ;
        RECT 31.265 17.135 31.515 20.665 ;
  LAYER M1 ;
        RECT 31.265 15.875 31.515 16.885 ;
  LAYER M1 ;
        RECT 31.265 11.255 31.515 14.785 ;
  LAYER M1 ;
        RECT 31.265 9.995 31.515 11.005 ;
  LAYER M1 ;
        RECT 31.265 7.895 31.515 8.905 ;
  LAYER M1 ;
        RECT 31.695 17.135 31.945 20.665 ;
  LAYER M1 ;
        RECT 31.695 11.255 31.945 14.785 ;
  LAYER M1 ;
        RECT 32.125 17.135 32.375 20.665 ;
  LAYER M1 ;
        RECT 32.125 15.875 32.375 16.885 ;
  LAYER M1 ;
        RECT 32.125 11.255 32.375 14.785 ;
  LAYER M1 ;
        RECT 32.125 9.995 32.375 11.005 ;
  LAYER M1 ;
        RECT 32.125 7.895 32.375 8.905 ;
  LAYER M1 ;
        RECT 32.555 17.135 32.805 20.665 ;
  LAYER M1 ;
        RECT 32.555 11.255 32.805 14.785 ;
  LAYER M1 ;
        RECT 32.985 17.135 33.235 20.665 ;
  LAYER M1 ;
        RECT 32.985 15.875 33.235 16.885 ;
  LAYER M1 ;
        RECT 32.985 11.255 33.235 14.785 ;
  LAYER M1 ;
        RECT 32.985 9.995 33.235 11.005 ;
  LAYER M1 ;
        RECT 32.985 7.895 33.235 8.905 ;
  LAYER M1 ;
        RECT 33.415 17.135 33.665 20.665 ;
  LAYER M1 ;
        RECT 33.415 11.255 33.665 14.785 ;
  LAYER M1 ;
        RECT 33.845 17.135 34.095 20.665 ;
  LAYER M1 ;
        RECT 33.845 15.875 34.095 16.885 ;
  LAYER M1 ;
        RECT 33.845 11.255 34.095 14.785 ;
  LAYER M1 ;
        RECT 33.845 9.995 34.095 11.005 ;
  LAYER M1 ;
        RECT 33.845 7.895 34.095 8.905 ;
  LAYER M1 ;
        RECT 34.275 17.135 34.525 20.665 ;
  LAYER M1 ;
        RECT 34.275 11.255 34.525 14.785 ;
  LAYER M1 ;
        RECT 34.705 17.135 34.955 20.665 ;
  LAYER M1 ;
        RECT 34.705 15.875 34.955 16.885 ;
  LAYER M1 ;
        RECT 34.705 11.255 34.955 14.785 ;
  LAYER M1 ;
        RECT 34.705 9.995 34.955 11.005 ;
  LAYER M1 ;
        RECT 34.705 7.895 34.955 8.905 ;
  LAYER M1 ;
        RECT 35.135 17.135 35.385 20.665 ;
  LAYER M1 ;
        RECT 35.135 11.255 35.385 14.785 ;
  LAYER M1 ;
        RECT 35.565 17.135 35.815 20.665 ;
  LAYER M1 ;
        RECT 35.565 15.875 35.815 16.885 ;
  LAYER M1 ;
        RECT 35.565 11.255 35.815 14.785 ;
  LAYER M1 ;
        RECT 35.565 9.995 35.815 11.005 ;
  LAYER M1 ;
        RECT 35.565 7.895 35.815 8.905 ;
  LAYER M1 ;
        RECT 35.995 17.135 36.245 20.665 ;
  LAYER M1 ;
        RECT 35.995 11.255 36.245 14.785 ;
  LAYER M2 ;
        RECT 26.06 20.44 35.86 20.72 ;
  LAYER M2 ;
        RECT 26.06 16.24 35.86 16.52 ;
  LAYER M2 ;
        RECT 25.63 20.02 36.29 20.3 ;
  LAYER M2 ;
        RECT 26.06 14.56 35.86 14.84 ;
  LAYER M2 ;
        RECT 26.06 10.36 35.86 10.64 ;
  LAYER M2 ;
        RECT 26.06 8.26 35.86 8.54 ;
  LAYER M2 ;
        RECT 25.63 14.14 36.29 14.42 ;
  LAYER M3 ;
        RECT 30.39 14.54 30.67 20.74 ;
  LAYER M3 ;
        RECT 30.82 10.34 31.1 16.54 ;
  LAYER M3 ;
        RECT 31.25 8.24 31.53 20.32 ;
  LAYER M1 ;
        RECT 11.485 17.135 11.735 20.665 ;
  LAYER M1 ;
        RECT 11.485 15.875 11.735 16.885 ;
  LAYER M1 ;
        RECT 11.485 11.255 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.485 9.995 11.735 11.005 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 8.905 ;
  LAYER M1 ;
        RECT 11.915 17.135 12.165 20.665 ;
  LAYER M1 ;
        RECT 11.915 11.255 12.165 14.785 ;
  LAYER M1 ;
        RECT 11.055 17.135 11.305 20.665 ;
  LAYER M1 ;
        RECT 11.055 11.255 11.305 14.785 ;
  LAYER M1 ;
        RECT 10.625 17.135 10.875 20.665 ;
  LAYER M1 ;
        RECT 10.625 15.875 10.875 16.885 ;
  LAYER M1 ;
        RECT 10.625 11.255 10.875 14.785 ;
  LAYER M1 ;
        RECT 10.625 9.995 10.875 11.005 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 8.905 ;
  LAYER M1 ;
        RECT 10.195 17.135 10.445 20.665 ;
  LAYER M1 ;
        RECT 10.195 11.255 10.445 14.785 ;
  LAYER M1 ;
        RECT 9.765 17.135 10.015 20.665 ;
  LAYER M1 ;
        RECT 9.765 15.875 10.015 16.885 ;
  LAYER M1 ;
        RECT 9.765 11.255 10.015 14.785 ;
  LAYER M1 ;
        RECT 9.765 9.995 10.015 11.005 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 8.905 ;
  LAYER M1 ;
        RECT 9.335 17.135 9.585 20.665 ;
  LAYER M1 ;
        RECT 9.335 11.255 9.585 14.785 ;
  LAYER M1 ;
        RECT 8.905 17.135 9.155 20.665 ;
  LAYER M1 ;
        RECT 8.905 15.875 9.155 16.885 ;
  LAYER M1 ;
        RECT 8.905 11.255 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.905 9.995 9.155 11.005 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 8.905 ;
  LAYER M1 ;
        RECT 8.475 17.135 8.725 20.665 ;
  LAYER M1 ;
        RECT 8.475 11.255 8.725 14.785 ;
  LAYER M1 ;
        RECT 8.045 17.135 8.295 20.665 ;
  LAYER M1 ;
        RECT 8.045 15.875 8.295 16.885 ;
  LAYER M1 ;
        RECT 8.045 11.255 8.295 14.785 ;
  LAYER M1 ;
        RECT 8.045 9.995 8.295 11.005 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 8.905 ;
  LAYER M1 ;
        RECT 7.615 17.135 7.865 20.665 ;
  LAYER M1 ;
        RECT 7.615 11.255 7.865 14.785 ;
  LAYER M1 ;
        RECT 7.185 17.135 7.435 20.665 ;
  LAYER M1 ;
        RECT 7.185 15.875 7.435 16.885 ;
  LAYER M1 ;
        RECT 7.185 11.255 7.435 14.785 ;
  LAYER M1 ;
        RECT 7.185 9.995 7.435 11.005 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.905 ;
  LAYER M1 ;
        RECT 6.755 17.135 7.005 20.665 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 6.325 17.135 6.575 20.665 ;
  LAYER M1 ;
        RECT 6.325 15.875 6.575 16.885 ;
  LAYER M1 ;
        RECT 6.325 11.255 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 11.005 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 8.905 ;
  LAYER M1 ;
        RECT 5.895 17.135 6.145 20.665 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M1 ;
        RECT 5.465 17.135 5.715 20.665 ;
  LAYER M1 ;
        RECT 5.465 15.875 5.715 16.885 ;
  LAYER M1 ;
        RECT 5.465 11.255 5.715 14.785 ;
  LAYER M1 ;
        RECT 5.465 9.995 5.715 11.005 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 8.905 ;
  LAYER M1 ;
        RECT 5.035 17.135 5.285 20.665 ;
  LAYER M1 ;
        RECT 5.035 11.255 5.285 14.785 ;
  LAYER M1 ;
        RECT 4.605 17.135 4.855 20.665 ;
  LAYER M1 ;
        RECT 4.605 15.875 4.855 16.885 ;
  LAYER M1 ;
        RECT 4.605 11.255 4.855 14.785 ;
  LAYER M1 ;
        RECT 4.605 9.995 4.855 11.005 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.905 ;
  LAYER M1 ;
        RECT 4.175 17.135 4.425 20.665 ;
  LAYER M1 ;
        RECT 4.175 11.255 4.425 14.785 ;
  LAYER M1 ;
        RECT 3.745 17.135 3.995 20.665 ;
  LAYER M1 ;
        RECT 3.745 15.875 3.995 16.885 ;
  LAYER M1 ;
        RECT 3.745 11.255 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.745 9.995 3.995 11.005 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 8.905 ;
  LAYER M1 ;
        RECT 3.315 17.135 3.565 20.665 ;
  LAYER M1 ;
        RECT 3.315 11.255 3.565 14.785 ;
  LAYER M1 ;
        RECT 2.885 17.135 3.135 20.665 ;
  LAYER M1 ;
        RECT 2.885 15.875 3.135 16.885 ;
  LAYER M1 ;
        RECT 2.885 11.255 3.135 14.785 ;
  LAYER M1 ;
        RECT 2.885 9.995 3.135 11.005 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.905 ;
  LAYER M1 ;
        RECT 2.455 17.135 2.705 20.665 ;
  LAYER M1 ;
        RECT 2.455 11.255 2.705 14.785 ;
  LAYER M1 ;
        RECT 2.025 17.135 2.275 20.665 ;
  LAYER M1 ;
        RECT 2.025 15.875 2.275 16.885 ;
  LAYER M1 ;
        RECT 2.025 11.255 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.025 9.995 2.275 11.005 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.905 ;
  LAYER M1 ;
        RECT 1.595 17.135 1.845 20.665 ;
  LAYER M1 ;
        RECT 1.595 11.255 1.845 14.785 ;
  LAYER M2 ;
        RECT 1.98 20.44 11.78 20.72 ;
  LAYER M2 ;
        RECT 1.98 16.24 11.78 16.52 ;
  LAYER M2 ;
        RECT 1.55 20.02 12.21 20.3 ;
  LAYER M2 ;
        RECT 1.98 14.56 11.78 14.84 ;
  LAYER M2 ;
        RECT 1.98 10.36 11.78 10.64 ;
  LAYER M2 ;
        RECT 1.98 8.26 11.78 8.54 ;
  LAYER M2 ;
        RECT 1.55 14.14 12.21 14.42 ;
  LAYER M3 ;
        RECT 7.17 14.54 7.45 20.74 ;
  LAYER M3 ;
        RECT 6.74 10.34 7.02 16.54 ;
  LAYER M3 ;
        RECT 6.31 8.24 6.59 20.32 ;
  LAYER M1 ;
        RECT 23.525 7.895 23.775 11.425 ;
  LAYER M1 ;
        RECT 23.525 11.675 23.775 12.685 ;
  LAYER M1 ;
        RECT 23.525 13.775 23.775 17.305 ;
  LAYER M1 ;
        RECT 23.525 17.555 23.775 18.565 ;
  LAYER M1 ;
        RECT 23.525 19.655 23.775 20.665 ;
  LAYER M1 ;
        RECT 23.955 7.895 24.205 11.425 ;
  LAYER M1 ;
        RECT 23.955 13.775 24.205 17.305 ;
  LAYER M1 ;
        RECT 23.095 7.895 23.345 11.425 ;
  LAYER M1 ;
        RECT 23.095 13.775 23.345 17.305 ;
  LAYER M1 ;
        RECT 22.665 7.895 22.915 11.425 ;
  LAYER M1 ;
        RECT 22.665 11.675 22.915 12.685 ;
  LAYER M1 ;
        RECT 22.665 13.775 22.915 17.305 ;
  LAYER M1 ;
        RECT 22.665 17.555 22.915 18.565 ;
  LAYER M1 ;
        RECT 22.665 19.655 22.915 20.665 ;
  LAYER M1 ;
        RECT 22.235 7.895 22.485 11.425 ;
  LAYER M1 ;
        RECT 22.235 13.775 22.485 17.305 ;
  LAYER M1 ;
        RECT 21.805 7.895 22.055 11.425 ;
  LAYER M1 ;
        RECT 21.805 11.675 22.055 12.685 ;
  LAYER M1 ;
        RECT 21.805 13.775 22.055 17.305 ;
  LAYER M1 ;
        RECT 21.805 17.555 22.055 18.565 ;
  LAYER M1 ;
        RECT 21.805 19.655 22.055 20.665 ;
  LAYER M1 ;
        RECT 21.375 7.895 21.625 11.425 ;
  LAYER M1 ;
        RECT 21.375 13.775 21.625 17.305 ;
  LAYER M1 ;
        RECT 20.945 7.895 21.195 11.425 ;
  LAYER M1 ;
        RECT 20.945 11.675 21.195 12.685 ;
  LAYER M1 ;
        RECT 20.945 13.775 21.195 17.305 ;
  LAYER M1 ;
        RECT 20.945 17.555 21.195 18.565 ;
  LAYER M1 ;
        RECT 20.945 19.655 21.195 20.665 ;
  LAYER M1 ;
        RECT 20.515 7.895 20.765 11.425 ;
  LAYER M1 ;
        RECT 20.515 13.775 20.765 17.305 ;
  LAYER M1 ;
        RECT 20.085 7.895 20.335 11.425 ;
  LAYER M1 ;
        RECT 20.085 11.675 20.335 12.685 ;
  LAYER M1 ;
        RECT 20.085 13.775 20.335 17.305 ;
  LAYER M1 ;
        RECT 20.085 17.555 20.335 18.565 ;
  LAYER M1 ;
        RECT 20.085 19.655 20.335 20.665 ;
  LAYER M1 ;
        RECT 19.655 7.895 19.905 11.425 ;
  LAYER M1 ;
        RECT 19.655 13.775 19.905 17.305 ;
  LAYER M2 ;
        RECT 20.04 7.84 23.82 8.12 ;
  LAYER M2 ;
        RECT 20.04 12.04 23.82 12.32 ;
  LAYER M2 ;
        RECT 19.61 8.26 24.25 8.54 ;
  LAYER M2 ;
        RECT 20.04 13.72 23.82 14 ;
  LAYER M2 ;
        RECT 20.04 17.92 23.82 18.2 ;
  LAYER M2 ;
        RECT 19.61 14.14 24.25 14.42 ;
  LAYER M2 ;
        RECT 20.04 20.02 23.82 20.3 ;
  LAYER M3 ;
        RECT 22.22 7.82 22.5 14.02 ;
  LAYER M3 ;
        RECT 21.79 12.02 22.07 18.22 ;
  LAYER M3 ;
        RECT 21.36 8.24 21.64 14.44 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 17.305 ;
  LAYER M1 ;
        RECT 14.065 17.555 14.315 18.565 ;
  LAYER M1 ;
        RECT 14.065 19.655 14.315 20.665 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 13.635 13.775 13.885 17.305 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M1 ;
        RECT 14.495 13.775 14.745 17.305 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 11.425 ;
  LAYER M1 ;
        RECT 14.925 11.675 15.175 12.685 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 17.305 ;
  LAYER M1 ;
        RECT 14.925 17.555 15.175 18.565 ;
  LAYER M1 ;
        RECT 14.925 19.655 15.175 20.665 ;
  LAYER M1 ;
        RECT 15.355 7.895 15.605 11.425 ;
  LAYER M1 ;
        RECT 15.355 13.775 15.605 17.305 ;
  LAYER M1 ;
        RECT 15.785 7.895 16.035 11.425 ;
  LAYER M1 ;
        RECT 15.785 11.675 16.035 12.685 ;
  LAYER M1 ;
        RECT 15.785 13.775 16.035 17.305 ;
  LAYER M1 ;
        RECT 15.785 17.555 16.035 18.565 ;
  LAYER M1 ;
        RECT 15.785 19.655 16.035 20.665 ;
  LAYER M1 ;
        RECT 16.215 7.895 16.465 11.425 ;
  LAYER M1 ;
        RECT 16.215 13.775 16.465 17.305 ;
  LAYER M1 ;
        RECT 16.645 7.895 16.895 11.425 ;
  LAYER M1 ;
        RECT 16.645 11.675 16.895 12.685 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 17.305 ;
  LAYER M1 ;
        RECT 16.645 17.555 16.895 18.565 ;
  LAYER M1 ;
        RECT 16.645 19.655 16.895 20.665 ;
  LAYER M1 ;
        RECT 17.075 7.895 17.325 11.425 ;
  LAYER M1 ;
        RECT 17.075 13.775 17.325 17.305 ;
  LAYER M1 ;
        RECT 17.505 7.895 17.755 11.425 ;
  LAYER M1 ;
        RECT 17.505 11.675 17.755 12.685 ;
  LAYER M1 ;
        RECT 17.505 13.775 17.755 17.305 ;
  LAYER M1 ;
        RECT 17.505 17.555 17.755 18.565 ;
  LAYER M1 ;
        RECT 17.505 19.655 17.755 20.665 ;
  LAYER M1 ;
        RECT 17.935 7.895 18.185 11.425 ;
  LAYER M1 ;
        RECT 17.935 13.775 18.185 17.305 ;
  LAYER M2 ;
        RECT 14.02 7.84 17.8 8.12 ;
  LAYER M2 ;
        RECT 14.02 12.04 17.8 12.32 ;
  LAYER M2 ;
        RECT 13.59 8.26 18.23 8.54 ;
  LAYER M2 ;
        RECT 14.02 13.72 17.8 14 ;
  LAYER M2 ;
        RECT 14.02 17.92 17.8 18.2 ;
  LAYER M2 ;
        RECT 13.59 14.14 18.23 14.42 ;
  LAYER M2 ;
        RECT 14.02 20.02 17.8 20.3 ;
  LAYER M3 ;
        RECT 15.34 7.82 15.62 14.02 ;
  LAYER M3 ;
        RECT 15.77 12.02 16.05 18.22 ;
  LAYER M3 ;
        RECT 16.2 8.24 16.48 14.44 ;
  END 
END CURRENT_MIRROR_OTA
