MACRO DCL_NMOS_S_42410075_X80_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_S_42410075_X80_Y1 0 0 ;
  SIZE 70520 BY 7560 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35120 260 35400 4780 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35550 680 35830 6880 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 7225 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 7225 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 7225 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 7225 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 7225 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 7225 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 7225 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8905 335 9155 3865 ;
    LAYER M1 ;
      RECT 8905 4115 9155 5125 ;
    LAYER M1 ;
      RECT 8905 6215 9155 7225 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 9765 335 10015 3865 ;
    LAYER M1 ;
      RECT 9765 4115 10015 5125 ;
    LAYER M1 ;
      RECT 9765 6215 10015 7225 ;
    LAYER M1 ;
      RECT 10195 335 10445 3865 ;
    LAYER M1 ;
      RECT 10625 335 10875 3865 ;
    LAYER M1 ;
      RECT 10625 4115 10875 5125 ;
    LAYER M1 ;
      RECT 10625 6215 10875 7225 ;
    LAYER M1 ;
      RECT 11055 335 11305 3865 ;
    LAYER M1 ;
      RECT 11485 335 11735 3865 ;
    LAYER M1 ;
      RECT 11485 4115 11735 5125 ;
    LAYER M1 ;
      RECT 11485 6215 11735 7225 ;
    LAYER M1 ;
      RECT 11915 335 12165 3865 ;
    LAYER M1 ;
      RECT 12345 335 12595 3865 ;
    LAYER M1 ;
      RECT 12345 4115 12595 5125 ;
    LAYER M1 ;
      RECT 12345 6215 12595 7225 ;
    LAYER M1 ;
      RECT 12775 335 13025 3865 ;
    LAYER M1 ;
      RECT 13205 335 13455 3865 ;
    LAYER M1 ;
      RECT 13205 4115 13455 5125 ;
    LAYER M1 ;
      RECT 13205 6215 13455 7225 ;
    LAYER M1 ;
      RECT 13635 335 13885 3865 ;
    LAYER M1 ;
      RECT 14065 335 14315 3865 ;
    LAYER M1 ;
      RECT 14065 4115 14315 5125 ;
    LAYER M1 ;
      RECT 14065 6215 14315 7225 ;
    LAYER M1 ;
      RECT 14495 335 14745 3865 ;
    LAYER M1 ;
      RECT 14925 335 15175 3865 ;
    LAYER M1 ;
      RECT 14925 4115 15175 5125 ;
    LAYER M1 ;
      RECT 14925 6215 15175 7225 ;
    LAYER M1 ;
      RECT 15355 335 15605 3865 ;
    LAYER M1 ;
      RECT 15785 335 16035 3865 ;
    LAYER M1 ;
      RECT 15785 4115 16035 5125 ;
    LAYER M1 ;
      RECT 15785 6215 16035 7225 ;
    LAYER M1 ;
      RECT 16215 335 16465 3865 ;
    LAYER M1 ;
      RECT 16645 335 16895 3865 ;
    LAYER M1 ;
      RECT 16645 4115 16895 5125 ;
    LAYER M1 ;
      RECT 16645 6215 16895 7225 ;
    LAYER M1 ;
      RECT 17075 335 17325 3865 ;
    LAYER M1 ;
      RECT 17505 335 17755 3865 ;
    LAYER M1 ;
      RECT 17505 4115 17755 5125 ;
    LAYER M1 ;
      RECT 17505 6215 17755 7225 ;
    LAYER M1 ;
      RECT 17935 335 18185 3865 ;
    LAYER M1 ;
      RECT 18365 335 18615 3865 ;
    LAYER M1 ;
      RECT 18365 4115 18615 5125 ;
    LAYER M1 ;
      RECT 18365 6215 18615 7225 ;
    LAYER M1 ;
      RECT 18795 335 19045 3865 ;
    LAYER M1 ;
      RECT 19225 335 19475 3865 ;
    LAYER M1 ;
      RECT 19225 4115 19475 5125 ;
    LAYER M1 ;
      RECT 19225 6215 19475 7225 ;
    LAYER M1 ;
      RECT 19655 335 19905 3865 ;
    LAYER M1 ;
      RECT 20085 335 20335 3865 ;
    LAYER M1 ;
      RECT 20085 4115 20335 5125 ;
    LAYER M1 ;
      RECT 20085 6215 20335 7225 ;
    LAYER M1 ;
      RECT 20515 335 20765 3865 ;
    LAYER M1 ;
      RECT 20945 335 21195 3865 ;
    LAYER M1 ;
      RECT 20945 4115 21195 5125 ;
    LAYER M1 ;
      RECT 20945 6215 21195 7225 ;
    LAYER M1 ;
      RECT 21375 335 21625 3865 ;
    LAYER M1 ;
      RECT 21805 335 22055 3865 ;
    LAYER M1 ;
      RECT 21805 4115 22055 5125 ;
    LAYER M1 ;
      RECT 21805 6215 22055 7225 ;
    LAYER M1 ;
      RECT 22235 335 22485 3865 ;
    LAYER M1 ;
      RECT 22665 335 22915 3865 ;
    LAYER M1 ;
      RECT 22665 4115 22915 5125 ;
    LAYER M1 ;
      RECT 22665 6215 22915 7225 ;
    LAYER M1 ;
      RECT 23095 335 23345 3865 ;
    LAYER M1 ;
      RECT 23525 335 23775 3865 ;
    LAYER M1 ;
      RECT 23525 4115 23775 5125 ;
    LAYER M1 ;
      RECT 23525 6215 23775 7225 ;
    LAYER M1 ;
      RECT 23955 335 24205 3865 ;
    LAYER M1 ;
      RECT 24385 335 24635 3865 ;
    LAYER M1 ;
      RECT 24385 4115 24635 5125 ;
    LAYER M1 ;
      RECT 24385 6215 24635 7225 ;
    LAYER M1 ;
      RECT 24815 335 25065 3865 ;
    LAYER M1 ;
      RECT 25245 335 25495 3865 ;
    LAYER M1 ;
      RECT 25245 4115 25495 5125 ;
    LAYER M1 ;
      RECT 25245 6215 25495 7225 ;
    LAYER M1 ;
      RECT 25675 335 25925 3865 ;
    LAYER M1 ;
      RECT 26105 335 26355 3865 ;
    LAYER M1 ;
      RECT 26105 4115 26355 5125 ;
    LAYER M1 ;
      RECT 26105 6215 26355 7225 ;
    LAYER M1 ;
      RECT 26535 335 26785 3865 ;
    LAYER M1 ;
      RECT 26965 335 27215 3865 ;
    LAYER M1 ;
      RECT 26965 4115 27215 5125 ;
    LAYER M1 ;
      RECT 26965 6215 27215 7225 ;
    LAYER M1 ;
      RECT 27395 335 27645 3865 ;
    LAYER M1 ;
      RECT 27825 335 28075 3865 ;
    LAYER M1 ;
      RECT 27825 4115 28075 5125 ;
    LAYER M1 ;
      RECT 27825 6215 28075 7225 ;
    LAYER M1 ;
      RECT 28255 335 28505 3865 ;
    LAYER M1 ;
      RECT 28685 335 28935 3865 ;
    LAYER M1 ;
      RECT 28685 4115 28935 5125 ;
    LAYER M1 ;
      RECT 28685 6215 28935 7225 ;
    LAYER M1 ;
      RECT 29115 335 29365 3865 ;
    LAYER M1 ;
      RECT 29545 335 29795 3865 ;
    LAYER M1 ;
      RECT 29545 4115 29795 5125 ;
    LAYER M1 ;
      RECT 29545 6215 29795 7225 ;
    LAYER M1 ;
      RECT 29975 335 30225 3865 ;
    LAYER M1 ;
      RECT 30405 335 30655 3865 ;
    LAYER M1 ;
      RECT 30405 4115 30655 5125 ;
    LAYER M1 ;
      RECT 30405 6215 30655 7225 ;
    LAYER M1 ;
      RECT 30835 335 31085 3865 ;
    LAYER M1 ;
      RECT 31265 335 31515 3865 ;
    LAYER M1 ;
      RECT 31265 4115 31515 5125 ;
    LAYER M1 ;
      RECT 31265 6215 31515 7225 ;
    LAYER M1 ;
      RECT 31695 335 31945 3865 ;
    LAYER M1 ;
      RECT 32125 335 32375 3865 ;
    LAYER M1 ;
      RECT 32125 4115 32375 5125 ;
    LAYER M1 ;
      RECT 32125 6215 32375 7225 ;
    LAYER M1 ;
      RECT 32555 335 32805 3865 ;
    LAYER M1 ;
      RECT 32985 335 33235 3865 ;
    LAYER M1 ;
      RECT 32985 4115 33235 5125 ;
    LAYER M1 ;
      RECT 32985 6215 33235 7225 ;
    LAYER M1 ;
      RECT 33415 335 33665 3865 ;
    LAYER M1 ;
      RECT 33845 335 34095 3865 ;
    LAYER M1 ;
      RECT 33845 4115 34095 5125 ;
    LAYER M1 ;
      RECT 33845 6215 34095 7225 ;
    LAYER M1 ;
      RECT 34275 335 34525 3865 ;
    LAYER M1 ;
      RECT 34705 335 34955 3865 ;
    LAYER M1 ;
      RECT 34705 4115 34955 5125 ;
    LAYER M1 ;
      RECT 34705 6215 34955 7225 ;
    LAYER M1 ;
      RECT 35135 335 35385 3865 ;
    LAYER M1 ;
      RECT 35565 335 35815 3865 ;
    LAYER M1 ;
      RECT 35565 4115 35815 5125 ;
    LAYER M1 ;
      RECT 35565 6215 35815 7225 ;
    LAYER M1 ;
      RECT 35995 335 36245 3865 ;
    LAYER M1 ;
      RECT 36425 335 36675 3865 ;
    LAYER M1 ;
      RECT 36425 4115 36675 5125 ;
    LAYER M1 ;
      RECT 36425 6215 36675 7225 ;
    LAYER M1 ;
      RECT 36855 335 37105 3865 ;
    LAYER M1 ;
      RECT 37285 335 37535 3865 ;
    LAYER M1 ;
      RECT 37285 4115 37535 5125 ;
    LAYER M1 ;
      RECT 37285 6215 37535 7225 ;
    LAYER M1 ;
      RECT 37715 335 37965 3865 ;
    LAYER M1 ;
      RECT 38145 335 38395 3865 ;
    LAYER M1 ;
      RECT 38145 4115 38395 5125 ;
    LAYER M1 ;
      RECT 38145 6215 38395 7225 ;
    LAYER M1 ;
      RECT 38575 335 38825 3865 ;
    LAYER M1 ;
      RECT 39005 335 39255 3865 ;
    LAYER M1 ;
      RECT 39005 4115 39255 5125 ;
    LAYER M1 ;
      RECT 39005 6215 39255 7225 ;
    LAYER M1 ;
      RECT 39435 335 39685 3865 ;
    LAYER M1 ;
      RECT 39865 335 40115 3865 ;
    LAYER M1 ;
      RECT 39865 4115 40115 5125 ;
    LAYER M1 ;
      RECT 39865 6215 40115 7225 ;
    LAYER M1 ;
      RECT 40295 335 40545 3865 ;
    LAYER M1 ;
      RECT 40725 335 40975 3865 ;
    LAYER M1 ;
      RECT 40725 4115 40975 5125 ;
    LAYER M1 ;
      RECT 40725 6215 40975 7225 ;
    LAYER M1 ;
      RECT 41155 335 41405 3865 ;
    LAYER M1 ;
      RECT 41585 335 41835 3865 ;
    LAYER M1 ;
      RECT 41585 4115 41835 5125 ;
    LAYER M1 ;
      RECT 41585 6215 41835 7225 ;
    LAYER M1 ;
      RECT 42015 335 42265 3865 ;
    LAYER M1 ;
      RECT 42445 335 42695 3865 ;
    LAYER M1 ;
      RECT 42445 4115 42695 5125 ;
    LAYER M1 ;
      RECT 42445 6215 42695 7225 ;
    LAYER M1 ;
      RECT 42875 335 43125 3865 ;
    LAYER M1 ;
      RECT 43305 335 43555 3865 ;
    LAYER M1 ;
      RECT 43305 4115 43555 5125 ;
    LAYER M1 ;
      RECT 43305 6215 43555 7225 ;
    LAYER M1 ;
      RECT 43735 335 43985 3865 ;
    LAYER M1 ;
      RECT 44165 335 44415 3865 ;
    LAYER M1 ;
      RECT 44165 4115 44415 5125 ;
    LAYER M1 ;
      RECT 44165 6215 44415 7225 ;
    LAYER M1 ;
      RECT 44595 335 44845 3865 ;
    LAYER M1 ;
      RECT 45025 335 45275 3865 ;
    LAYER M1 ;
      RECT 45025 4115 45275 5125 ;
    LAYER M1 ;
      RECT 45025 6215 45275 7225 ;
    LAYER M1 ;
      RECT 45455 335 45705 3865 ;
    LAYER M1 ;
      RECT 45885 335 46135 3865 ;
    LAYER M1 ;
      RECT 45885 4115 46135 5125 ;
    LAYER M1 ;
      RECT 45885 6215 46135 7225 ;
    LAYER M1 ;
      RECT 46315 335 46565 3865 ;
    LAYER M1 ;
      RECT 46745 335 46995 3865 ;
    LAYER M1 ;
      RECT 46745 4115 46995 5125 ;
    LAYER M1 ;
      RECT 46745 6215 46995 7225 ;
    LAYER M1 ;
      RECT 47175 335 47425 3865 ;
    LAYER M1 ;
      RECT 47605 335 47855 3865 ;
    LAYER M1 ;
      RECT 47605 4115 47855 5125 ;
    LAYER M1 ;
      RECT 47605 6215 47855 7225 ;
    LAYER M1 ;
      RECT 48035 335 48285 3865 ;
    LAYER M1 ;
      RECT 48465 335 48715 3865 ;
    LAYER M1 ;
      RECT 48465 4115 48715 5125 ;
    LAYER M1 ;
      RECT 48465 6215 48715 7225 ;
    LAYER M1 ;
      RECT 48895 335 49145 3865 ;
    LAYER M1 ;
      RECT 49325 335 49575 3865 ;
    LAYER M1 ;
      RECT 49325 4115 49575 5125 ;
    LAYER M1 ;
      RECT 49325 6215 49575 7225 ;
    LAYER M1 ;
      RECT 49755 335 50005 3865 ;
    LAYER M1 ;
      RECT 50185 335 50435 3865 ;
    LAYER M1 ;
      RECT 50185 4115 50435 5125 ;
    LAYER M1 ;
      RECT 50185 6215 50435 7225 ;
    LAYER M1 ;
      RECT 50615 335 50865 3865 ;
    LAYER M1 ;
      RECT 51045 335 51295 3865 ;
    LAYER M1 ;
      RECT 51045 4115 51295 5125 ;
    LAYER M1 ;
      RECT 51045 6215 51295 7225 ;
    LAYER M1 ;
      RECT 51475 335 51725 3865 ;
    LAYER M1 ;
      RECT 51905 335 52155 3865 ;
    LAYER M1 ;
      RECT 51905 4115 52155 5125 ;
    LAYER M1 ;
      RECT 51905 6215 52155 7225 ;
    LAYER M1 ;
      RECT 52335 335 52585 3865 ;
    LAYER M1 ;
      RECT 52765 335 53015 3865 ;
    LAYER M1 ;
      RECT 52765 4115 53015 5125 ;
    LAYER M1 ;
      RECT 52765 6215 53015 7225 ;
    LAYER M1 ;
      RECT 53195 335 53445 3865 ;
    LAYER M1 ;
      RECT 53625 335 53875 3865 ;
    LAYER M1 ;
      RECT 53625 4115 53875 5125 ;
    LAYER M1 ;
      RECT 53625 6215 53875 7225 ;
    LAYER M1 ;
      RECT 54055 335 54305 3865 ;
    LAYER M1 ;
      RECT 54485 335 54735 3865 ;
    LAYER M1 ;
      RECT 54485 4115 54735 5125 ;
    LAYER M1 ;
      RECT 54485 6215 54735 7225 ;
    LAYER M1 ;
      RECT 54915 335 55165 3865 ;
    LAYER M1 ;
      RECT 55345 335 55595 3865 ;
    LAYER M1 ;
      RECT 55345 4115 55595 5125 ;
    LAYER M1 ;
      RECT 55345 6215 55595 7225 ;
    LAYER M1 ;
      RECT 55775 335 56025 3865 ;
    LAYER M1 ;
      RECT 56205 335 56455 3865 ;
    LAYER M1 ;
      RECT 56205 4115 56455 5125 ;
    LAYER M1 ;
      RECT 56205 6215 56455 7225 ;
    LAYER M1 ;
      RECT 56635 335 56885 3865 ;
    LAYER M1 ;
      RECT 57065 335 57315 3865 ;
    LAYER M1 ;
      RECT 57065 4115 57315 5125 ;
    LAYER M1 ;
      RECT 57065 6215 57315 7225 ;
    LAYER M1 ;
      RECT 57495 335 57745 3865 ;
    LAYER M1 ;
      RECT 57925 335 58175 3865 ;
    LAYER M1 ;
      RECT 57925 4115 58175 5125 ;
    LAYER M1 ;
      RECT 57925 6215 58175 7225 ;
    LAYER M1 ;
      RECT 58355 335 58605 3865 ;
    LAYER M1 ;
      RECT 58785 335 59035 3865 ;
    LAYER M1 ;
      RECT 58785 4115 59035 5125 ;
    LAYER M1 ;
      RECT 58785 6215 59035 7225 ;
    LAYER M1 ;
      RECT 59215 335 59465 3865 ;
    LAYER M1 ;
      RECT 59645 335 59895 3865 ;
    LAYER M1 ;
      RECT 59645 4115 59895 5125 ;
    LAYER M1 ;
      RECT 59645 6215 59895 7225 ;
    LAYER M1 ;
      RECT 60075 335 60325 3865 ;
    LAYER M1 ;
      RECT 60505 335 60755 3865 ;
    LAYER M1 ;
      RECT 60505 4115 60755 5125 ;
    LAYER M1 ;
      RECT 60505 6215 60755 7225 ;
    LAYER M1 ;
      RECT 60935 335 61185 3865 ;
    LAYER M1 ;
      RECT 61365 335 61615 3865 ;
    LAYER M1 ;
      RECT 61365 4115 61615 5125 ;
    LAYER M1 ;
      RECT 61365 6215 61615 7225 ;
    LAYER M1 ;
      RECT 61795 335 62045 3865 ;
    LAYER M1 ;
      RECT 62225 335 62475 3865 ;
    LAYER M1 ;
      RECT 62225 4115 62475 5125 ;
    LAYER M1 ;
      RECT 62225 6215 62475 7225 ;
    LAYER M1 ;
      RECT 62655 335 62905 3865 ;
    LAYER M1 ;
      RECT 63085 335 63335 3865 ;
    LAYER M1 ;
      RECT 63085 4115 63335 5125 ;
    LAYER M1 ;
      RECT 63085 6215 63335 7225 ;
    LAYER M1 ;
      RECT 63515 335 63765 3865 ;
    LAYER M1 ;
      RECT 63945 335 64195 3865 ;
    LAYER M1 ;
      RECT 63945 4115 64195 5125 ;
    LAYER M1 ;
      RECT 63945 6215 64195 7225 ;
    LAYER M1 ;
      RECT 64375 335 64625 3865 ;
    LAYER M1 ;
      RECT 64805 335 65055 3865 ;
    LAYER M1 ;
      RECT 64805 4115 65055 5125 ;
    LAYER M1 ;
      RECT 64805 6215 65055 7225 ;
    LAYER M1 ;
      RECT 65235 335 65485 3865 ;
    LAYER M1 ;
      RECT 65665 335 65915 3865 ;
    LAYER M1 ;
      RECT 65665 4115 65915 5125 ;
    LAYER M1 ;
      RECT 65665 6215 65915 7225 ;
    LAYER M1 ;
      RECT 66095 335 66345 3865 ;
    LAYER M1 ;
      RECT 66525 335 66775 3865 ;
    LAYER M1 ;
      RECT 66525 4115 66775 5125 ;
    LAYER M1 ;
      RECT 66525 6215 66775 7225 ;
    LAYER M1 ;
      RECT 66955 335 67205 3865 ;
    LAYER M1 ;
      RECT 67385 335 67635 3865 ;
    LAYER M1 ;
      RECT 67385 4115 67635 5125 ;
    LAYER M1 ;
      RECT 67385 6215 67635 7225 ;
    LAYER M1 ;
      RECT 67815 335 68065 3865 ;
    LAYER M1 ;
      RECT 68245 335 68495 3865 ;
    LAYER M1 ;
      RECT 68245 4115 68495 5125 ;
    LAYER M1 ;
      RECT 68245 6215 68495 7225 ;
    LAYER M1 ;
      RECT 68675 335 68925 3865 ;
    LAYER M1 ;
      RECT 69105 335 69355 3865 ;
    LAYER M1 ;
      RECT 69105 4115 69355 5125 ;
    LAYER M1 ;
      RECT 69105 6215 69355 7225 ;
    LAYER M1 ;
      RECT 69535 335 69785 3865 ;
    LAYER M2 ;
      RECT 1120 4480 69400 4760 ;
    LAYER M2 ;
      RECT 1120 280 69400 560 ;
    LAYER M2 ;
      RECT 1120 6580 69400 6860 ;
    LAYER M2 ;
      RECT 690 700 69830 980 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6635 3095 6805 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6635 3955 6805 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6635 4815 6805 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6635 5675 6805 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6635 6535 6805 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6635 7395 6805 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6635 8255 6805 ;
    LAYER V1 ;
      RECT 8945 335 9115 505 ;
    LAYER V1 ;
      RECT 8945 4535 9115 4705 ;
    LAYER V1 ;
      RECT 8945 6635 9115 6805 ;
    LAYER V1 ;
      RECT 9805 335 9975 505 ;
    LAYER V1 ;
      RECT 9805 4535 9975 4705 ;
    LAYER V1 ;
      RECT 9805 6635 9975 6805 ;
    LAYER V1 ;
      RECT 10665 335 10835 505 ;
    LAYER V1 ;
      RECT 10665 4535 10835 4705 ;
    LAYER V1 ;
      RECT 10665 6635 10835 6805 ;
    LAYER V1 ;
      RECT 11525 335 11695 505 ;
    LAYER V1 ;
      RECT 11525 4535 11695 4705 ;
    LAYER V1 ;
      RECT 11525 6635 11695 6805 ;
    LAYER V1 ;
      RECT 12385 335 12555 505 ;
    LAYER V1 ;
      RECT 12385 4535 12555 4705 ;
    LAYER V1 ;
      RECT 12385 6635 12555 6805 ;
    LAYER V1 ;
      RECT 13245 335 13415 505 ;
    LAYER V1 ;
      RECT 13245 4535 13415 4705 ;
    LAYER V1 ;
      RECT 13245 6635 13415 6805 ;
    LAYER V1 ;
      RECT 14105 335 14275 505 ;
    LAYER V1 ;
      RECT 14105 4535 14275 4705 ;
    LAYER V1 ;
      RECT 14105 6635 14275 6805 ;
    LAYER V1 ;
      RECT 14965 335 15135 505 ;
    LAYER V1 ;
      RECT 14965 4535 15135 4705 ;
    LAYER V1 ;
      RECT 14965 6635 15135 6805 ;
    LAYER V1 ;
      RECT 15825 335 15995 505 ;
    LAYER V1 ;
      RECT 15825 4535 15995 4705 ;
    LAYER V1 ;
      RECT 15825 6635 15995 6805 ;
    LAYER V1 ;
      RECT 16685 335 16855 505 ;
    LAYER V1 ;
      RECT 16685 4535 16855 4705 ;
    LAYER V1 ;
      RECT 16685 6635 16855 6805 ;
    LAYER V1 ;
      RECT 17545 335 17715 505 ;
    LAYER V1 ;
      RECT 17545 4535 17715 4705 ;
    LAYER V1 ;
      RECT 17545 6635 17715 6805 ;
    LAYER V1 ;
      RECT 18405 335 18575 505 ;
    LAYER V1 ;
      RECT 18405 4535 18575 4705 ;
    LAYER V1 ;
      RECT 18405 6635 18575 6805 ;
    LAYER V1 ;
      RECT 19265 335 19435 505 ;
    LAYER V1 ;
      RECT 19265 4535 19435 4705 ;
    LAYER V1 ;
      RECT 19265 6635 19435 6805 ;
    LAYER V1 ;
      RECT 20125 335 20295 505 ;
    LAYER V1 ;
      RECT 20125 4535 20295 4705 ;
    LAYER V1 ;
      RECT 20125 6635 20295 6805 ;
    LAYER V1 ;
      RECT 20985 335 21155 505 ;
    LAYER V1 ;
      RECT 20985 4535 21155 4705 ;
    LAYER V1 ;
      RECT 20985 6635 21155 6805 ;
    LAYER V1 ;
      RECT 21845 335 22015 505 ;
    LAYER V1 ;
      RECT 21845 4535 22015 4705 ;
    LAYER V1 ;
      RECT 21845 6635 22015 6805 ;
    LAYER V1 ;
      RECT 22705 335 22875 505 ;
    LAYER V1 ;
      RECT 22705 4535 22875 4705 ;
    LAYER V1 ;
      RECT 22705 6635 22875 6805 ;
    LAYER V1 ;
      RECT 23565 335 23735 505 ;
    LAYER V1 ;
      RECT 23565 4535 23735 4705 ;
    LAYER V1 ;
      RECT 23565 6635 23735 6805 ;
    LAYER V1 ;
      RECT 24425 335 24595 505 ;
    LAYER V1 ;
      RECT 24425 4535 24595 4705 ;
    LAYER V1 ;
      RECT 24425 6635 24595 6805 ;
    LAYER V1 ;
      RECT 25285 335 25455 505 ;
    LAYER V1 ;
      RECT 25285 4535 25455 4705 ;
    LAYER V1 ;
      RECT 25285 6635 25455 6805 ;
    LAYER V1 ;
      RECT 26145 335 26315 505 ;
    LAYER V1 ;
      RECT 26145 4535 26315 4705 ;
    LAYER V1 ;
      RECT 26145 6635 26315 6805 ;
    LAYER V1 ;
      RECT 27005 335 27175 505 ;
    LAYER V1 ;
      RECT 27005 4535 27175 4705 ;
    LAYER V1 ;
      RECT 27005 6635 27175 6805 ;
    LAYER V1 ;
      RECT 27865 335 28035 505 ;
    LAYER V1 ;
      RECT 27865 4535 28035 4705 ;
    LAYER V1 ;
      RECT 27865 6635 28035 6805 ;
    LAYER V1 ;
      RECT 28725 335 28895 505 ;
    LAYER V1 ;
      RECT 28725 4535 28895 4705 ;
    LAYER V1 ;
      RECT 28725 6635 28895 6805 ;
    LAYER V1 ;
      RECT 29585 335 29755 505 ;
    LAYER V1 ;
      RECT 29585 4535 29755 4705 ;
    LAYER V1 ;
      RECT 29585 6635 29755 6805 ;
    LAYER V1 ;
      RECT 30445 335 30615 505 ;
    LAYER V1 ;
      RECT 30445 4535 30615 4705 ;
    LAYER V1 ;
      RECT 30445 6635 30615 6805 ;
    LAYER V1 ;
      RECT 31305 335 31475 505 ;
    LAYER V1 ;
      RECT 31305 4535 31475 4705 ;
    LAYER V1 ;
      RECT 31305 6635 31475 6805 ;
    LAYER V1 ;
      RECT 32165 335 32335 505 ;
    LAYER V1 ;
      RECT 32165 4535 32335 4705 ;
    LAYER V1 ;
      RECT 32165 6635 32335 6805 ;
    LAYER V1 ;
      RECT 33025 335 33195 505 ;
    LAYER V1 ;
      RECT 33025 4535 33195 4705 ;
    LAYER V1 ;
      RECT 33025 6635 33195 6805 ;
    LAYER V1 ;
      RECT 33885 335 34055 505 ;
    LAYER V1 ;
      RECT 33885 4535 34055 4705 ;
    LAYER V1 ;
      RECT 33885 6635 34055 6805 ;
    LAYER V1 ;
      RECT 34745 335 34915 505 ;
    LAYER V1 ;
      RECT 34745 4535 34915 4705 ;
    LAYER V1 ;
      RECT 34745 6635 34915 6805 ;
    LAYER V1 ;
      RECT 35605 335 35775 505 ;
    LAYER V1 ;
      RECT 35605 4535 35775 4705 ;
    LAYER V1 ;
      RECT 35605 6635 35775 6805 ;
    LAYER V1 ;
      RECT 36465 335 36635 505 ;
    LAYER V1 ;
      RECT 36465 4535 36635 4705 ;
    LAYER V1 ;
      RECT 36465 6635 36635 6805 ;
    LAYER V1 ;
      RECT 37325 335 37495 505 ;
    LAYER V1 ;
      RECT 37325 4535 37495 4705 ;
    LAYER V1 ;
      RECT 37325 6635 37495 6805 ;
    LAYER V1 ;
      RECT 38185 335 38355 505 ;
    LAYER V1 ;
      RECT 38185 4535 38355 4705 ;
    LAYER V1 ;
      RECT 38185 6635 38355 6805 ;
    LAYER V1 ;
      RECT 39045 335 39215 505 ;
    LAYER V1 ;
      RECT 39045 4535 39215 4705 ;
    LAYER V1 ;
      RECT 39045 6635 39215 6805 ;
    LAYER V1 ;
      RECT 39905 335 40075 505 ;
    LAYER V1 ;
      RECT 39905 4535 40075 4705 ;
    LAYER V1 ;
      RECT 39905 6635 40075 6805 ;
    LAYER V1 ;
      RECT 40765 335 40935 505 ;
    LAYER V1 ;
      RECT 40765 4535 40935 4705 ;
    LAYER V1 ;
      RECT 40765 6635 40935 6805 ;
    LAYER V1 ;
      RECT 41625 335 41795 505 ;
    LAYER V1 ;
      RECT 41625 4535 41795 4705 ;
    LAYER V1 ;
      RECT 41625 6635 41795 6805 ;
    LAYER V1 ;
      RECT 42485 335 42655 505 ;
    LAYER V1 ;
      RECT 42485 4535 42655 4705 ;
    LAYER V1 ;
      RECT 42485 6635 42655 6805 ;
    LAYER V1 ;
      RECT 43345 335 43515 505 ;
    LAYER V1 ;
      RECT 43345 4535 43515 4705 ;
    LAYER V1 ;
      RECT 43345 6635 43515 6805 ;
    LAYER V1 ;
      RECT 44205 335 44375 505 ;
    LAYER V1 ;
      RECT 44205 4535 44375 4705 ;
    LAYER V1 ;
      RECT 44205 6635 44375 6805 ;
    LAYER V1 ;
      RECT 45065 335 45235 505 ;
    LAYER V1 ;
      RECT 45065 4535 45235 4705 ;
    LAYER V1 ;
      RECT 45065 6635 45235 6805 ;
    LAYER V1 ;
      RECT 45925 335 46095 505 ;
    LAYER V1 ;
      RECT 45925 4535 46095 4705 ;
    LAYER V1 ;
      RECT 45925 6635 46095 6805 ;
    LAYER V1 ;
      RECT 46785 335 46955 505 ;
    LAYER V1 ;
      RECT 46785 4535 46955 4705 ;
    LAYER V1 ;
      RECT 46785 6635 46955 6805 ;
    LAYER V1 ;
      RECT 47645 335 47815 505 ;
    LAYER V1 ;
      RECT 47645 4535 47815 4705 ;
    LAYER V1 ;
      RECT 47645 6635 47815 6805 ;
    LAYER V1 ;
      RECT 48505 335 48675 505 ;
    LAYER V1 ;
      RECT 48505 4535 48675 4705 ;
    LAYER V1 ;
      RECT 48505 6635 48675 6805 ;
    LAYER V1 ;
      RECT 49365 335 49535 505 ;
    LAYER V1 ;
      RECT 49365 4535 49535 4705 ;
    LAYER V1 ;
      RECT 49365 6635 49535 6805 ;
    LAYER V1 ;
      RECT 50225 335 50395 505 ;
    LAYER V1 ;
      RECT 50225 4535 50395 4705 ;
    LAYER V1 ;
      RECT 50225 6635 50395 6805 ;
    LAYER V1 ;
      RECT 51085 335 51255 505 ;
    LAYER V1 ;
      RECT 51085 4535 51255 4705 ;
    LAYER V1 ;
      RECT 51085 6635 51255 6805 ;
    LAYER V1 ;
      RECT 51945 335 52115 505 ;
    LAYER V1 ;
      RECT 51945 4535 52115 4705 ;
    LAYER V1 ;
      RECT 51945 6635 52115 6805 ;
    LAYER V1 ;
      RECT 52805 335 52975 505 ;
    LAYER V1 ;
      RECT 52805 4535 52975 4705 ;
    LAYER V1 ;
      RECT 52805 6635 52975 6805 ;
    LAYER V1 ;
      RECT 53665 335 53835 505 ;
    LAYER V1 ;
      RECT 53665 4535 53835 4705 ;
    LAYER V1 ;
      RECT 53665 6635 53835 6805 ;
    LAYER V1 ;
      RECT 54525 335 54695 505 ;
    LAYER V1 ;
      RECT 54525 4535 54695 4705 ;
    LAYER V1 ;
      RECT 54525 6635 54695 6805 ;
    LAYER V1 ;
      RECT 55385 335 55555 505 ;
    LAYER V1 ;
      RECT 55385 4535 55555 4705 ;
    LAYER V1 ;
      RECT 55385 6635 55555 6805 ;
    LAYER V1 ;
      RECT 56245 335 56415 505 ;
    LAYER V1 ;
      RECT 56245 4535 56415 4705 ;
    LAYER V1 ;
      RECT 56245 6635 56415 6805 ;
    LAYER V1 ;
      RECT 57105 335 57275 505 ;
    LAYER V1 ;
      RECT 57105 4535 57275 4705 ;
    LAYER V1 ;
      RECT 57105 6635 57275 6805 ;
    LAYER V1 ;
      RECT 57965 335 58135 505 ;
    LAYER V1 ;
      RECT 57965 4535 58135 4705 ;
    LAYER V1 ;
      RECT 57965 6635 58135 6805 ;
    LAYER V1 ;
      RECT 58825 335 58995 505 ;
    LAYER V1 ;
      RECT 58825 4535 58995 4705 ;
    LAYER V1 ;
      RECT 58825 6635 58995 6805 ;
    LAYER V1 ;
      RECT 59685 335 59855 505 ;
    LAYER V1 ;
      RECT 59685 4535 59855 4705 ;
    LAYER V1 ;
      RECT 59685 6635 59855 6805 ;
    LAYER V1 ;
      RECT 60545 335 60715 505 ;
    LAYER V1 ;
      RECT 60545 4535 60715 4705 ;
    LAYER V1 ;
      RECT 60545 6635 60715 6805 ;
    LAYER V1 ;
      RECT 61405 335 61575 505 ;
    LAYER V1 ;
      RECT 61405 4535 61575 4705 ;
    LAYER V1 ;
      RECT 61405 6635 61575 6805 ;
    LAYER V1 ;
      RECT 62265 335 62435 505 ;
    LAYER V1 ;
      RECT 62265 4535 62435 4705 ;
    LAYER V1 ;
      RECT 62265 6635 62435 6805 ;
    LAYER V1 ;
      RECT 63125 335 63295 505 ;
    LAYER V1 ;
      RECT 63125 4535 63295 4705 ;
    LAYER V1 ;
      RECT 63125 6635 63295 6805 ;
    LAYER V1 ;
      RECT 63985 335 64155 505 ;
    LAYER V1 ;
      RECT 63985 4535 64155 4705 ;
    LAYER V1 ;
      RECT 63985 6635 64155 6805 ;
    LAYER V1 ;
      RECT 64845 335 65015 505 ;
    LAYER V1 ;
      RECT 64845 4535 65015 4705 ;
    LAYER V1 ;
      RECT 64845 6635 65015 6805 ;
    LAYER V1 ;
      RECT 65705 335 65875 505 ;
    LAYER V1 ;
      RECT 65705 4535 65875 4705 ;
    LAYER V1 ;
      RECT 65705 6635 65875 6805 ;
    LAYER V1 ;
      RECT 66565 335 66735 505 ;
    LAYER V1 ;
      RECT 66565 4535 66735 4705 ;
    LAYER V1 ;
      RECT 66565 6635 66735 6805 ;
    LAYER V1 ;
      RECT 67425 335 67595 505 ;
    LAYER V1 ;
      RECT 67425 4535 67595 4705 ;
    LAYER V1 ;
      RECT 67425 6635 67595 6805 ;
    LAYER V1 ;
      RECT 68285 335 68455 505 ;
    LAYER V1 ;
      RECT 68285 4535 68455 4705 ;
    LAYER V1 ;
      RECT 68285 6635 68455 6805 ;
    LAYER V1 ;
      RECT 69145 335 69315 505 ;
    LAYER V1 ;
      RECT 69145 4535 69315 4705 ;
    LAYER V1 ;
      RECT 69145 6635 69315 6805 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 8515 755 8685 925 ;
    LAYER V1 ;
      RECT 9375 755 9545 925 ;
    LAYER V1 ;
      RECT 10235 755 10405 925 ;
    LAYER V1 ;
      RECT 11095 755 11265 925 ;
    LAYER V1 ;
      RECT 11955 755 12125 925 ;
    LAYER V1 ;
      RECT 12815 755 12985 925 ;
    LAYER V1 ;
      RECT 13675 755 13845 925 ;
    LAYER V1 ;
      RECT 14535 755 14705 925 ;
    LAYER V1 ;
      RECT 15395 755 15565 925 ;
    LAYER V1 ;
      RECT 16255 755 16425 925 ;
    LAYER V1 ;
      RECT 17115 755 17285 925 ;
    LAYER V1 ;
      RECT 17975 755 18145 925 ;
    LAYER V1 ;
      RECT 18835 755 19005 925 ;
    LAYER V1 ;
      RECT 19695 755 19865 925 ;
    LAYER V1 ;
      RECT 20555 755 20725 925 ;
    LAYER V1 ;
      RECT 21415 755 21585 925 ;
    LAYER V1 ;
      RECT 22275 755 22445 925 ;
    LAYER V1 ;
      RECT 23135 755 23305 925 ;
    LAYER V1 ;
      RECT 23995 755 24165 925 ;
    LAYER V1 ;
      RECT 24855 755 25025 925 ;
    LAYER V1 ;
      RECT 25715 755 25885 925 ;
    LAYER V1 ;
      RECT 26575 755 26745 925 ;
    LAYER V1 ;
      RECT 27435 755 27605 925 ;
    LAYER V1 ;
      RECT 28295 755 28465 925 ;
    LAYER V1 ;
      RECT 29155 755 29325 925 ;
    LAYER V1 ;
      RECT 30015 755 30185 925 ;
    LAYER V1 ;
      RECT 30875 755 31045 925 ;
    LAYER V1 ;
      RECT 31735 755 31905 925 ;
    LAYER V1 ;
      RECT 32595 755 32765 925 ;
    LAYER V1 ;
      RECT 33455 755 33625 925 ;
    LAYER V1 ;
      RECT 34315 755 34485 925 ;
    LAYER V1 ;
      RECT 35175 755 35345 925 ;
    LAYER V1 ;
      RECT 36035 755 36205 925 ;
    LAYER V1 ;
      RECT 36895 755 37065 925 ;
    LAYER V1 ;
      RECT 37755 755 37925 925 ;
    LAYER V1 ;
      RECT 38615 755 38785 925 ;
    LAYER V1 ;
      RECT 39475 755 39645 925 ;
    LAYER V1 ;
      RECT 40335 755 40505 925 ;
    LAYER V1 ;
      RECT 41195 755 41365 925 ;
    LAYER V1 ;
      RECT 42055 755 42225 925 ;
    LAYER V1 ;
      RECT 42915 755 43085 925 ;
    LAYER V1 ;
      RECT 43775 755 43945 925 ;
    LAYER V1 ;
      RECT 44635 755 44805 925 ;
    LAYER V1 ;
      RECT 45495 755 45665 925 ;
    LAYER V1 ;
      RECT 46355 755 46525 925 ;
    LAYER V1 ;
      RECT 47215 755 47385 925 ;
    LAYER V1 ;
      RECT 48075 755 48245 925 ;
    LAYER V1 ;
      RECT 48935 755 49105 925 ;
    LAYER V1 ;
      RECT 49795 755 49965 925 ;
    LAYER V1 ;
      RECT 50655 755 50825 925 ;
    LAYER V1 ;
      RECT 51515 755 51685 925 ;
    LAYER V1 ;
      RECT 52375 755 52545 925 ;
    LAYER V1 ;
      RECT 53235 755 53405 925 ;
    LAYER V1 ;
      RECT 54095 755 54265 925 ;
    LAYER V1 ;
      RECT 54955 755 55125 925 ;
    LAYER V1 ;
      RECT 55815 755 55985 925 ;
    LAYER V1 ;
      RECT 56675 755 56845 925 ;
    LAYER V1 ;
      RECT 57535 755 57705 925 ;
    LAYER V1 ;
      RECT 58395 755 58565 925 ;
    LAYER V1 ;
      RECT 59255 755 59425 925 ;
    LAYER V1 ;
      RECT 60115 755 60285 925 ;
    LAYER V1 ;
      RECT 60975 755 61145 925 ;
    LAYER V1 ;
      RECT 61835 755 62005 925 ;
    LAYER V1 ;
      RECT 62695 755 62865 925 ;
    LAYER V1 ;
      RECT 63555 755 63725 925 ;
    LAYER V1 ;
      RECT 64415 755 64585 925 ;
    LAYER V1 ;
      RECT 65275 755 65445 925 ;
    LAYER V1 ;
      RECT 66135 755 66305 925 ;
    LAYER V1 ;
      RECT 66995 755 67165 925 ;
    LAYER V1 ;
      RECT 67855 755 68025 925 ;
    LAYER V1 ;
      RECT 68715 755 68885 925 ;
    LAYER V1 ;
      RECT 69575 755 69745 925 ;
    LAYER V2 ;
      RECT 35185 345 35335 495 ;
    LAYER V2 ;
      RECT 35185 4545 35335 4695 ;
    LAYER V2 ;
      RECT 35615 765 35765 915 ;
    LAYER V2 ;
      RECT 35615 6645 35765 6795 ;
  END
END DCL_NMOS_S_42410075_X80_Y1
