MACRO DCL_NMOS_S_42410075_X2_Y40
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_S_42410075_X2_Y40 0 0 ;
  SIZE 3440 BY 236880 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 260 1860 234100 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 680 2290 236200 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 62665 ;
    LAYER M1 ;
      RECT 1165 62915 1415 63925 ;
    LAYER M1 ;
      RECT 1165 65015 1415 68545 ;
    LAYER M1 ;
      RECT 1165 68795 1415 69805 ;
    LAYER M1 ;
      RECT 1165 70895 1415 74425 ;
    LAYER M1 ;
      RECT 1165 74675 1415 75685 ;
    LAYER M1 ;
      RECT 1165 76775 1415 80305 ;
    LAYER M1 ;
      RECT 1165 80555 1415 81565 ;
    LAYER M1 ;
      RECT 1165 82655 1415 86185 ;
    LAYER M1 ;
      RECT 1165 86435 1415 87445 ;
    LAYER M1 ;
      RECT 1165 88535 1415 92065 ;
    LAYER M1 ;
      RECT 1165 92315 1415 93325 ;
    LAYER M1 ;
      RECT 1165 94415 1415 97945 ;
    LAYER M1 ;
      RECT 1165 98195 1415 99205 ;
    LAYER M1 ;
      RECT 1165 100295 1415 103825 ;
    LAYER M1 ;
      RECT 1165 104075 1415 105085 ;
    LAYER M1 ;
      RECT 1165 106175 1415 109705 ;
    LAYER M1 ;
      RECT 1165 109955 1415 110965 ;
    LAYER M1 ;
      RECT 1165 112055 1415 115585 ;
    LAYER M1 ;
      RECT 1165 115835 1415 116845 ;
    LAYER M1 ;
      RECT 1165 117935 1415 121465 ;
    LAYER M1 ;
      RECT 1165 121715 1415 122725 ;
    LAYER M1 ;
      RECT 1165 123815 1415 127345 ;
    LAYER M1 ;
      RECT 1165 127595 1415 128605 ;
    LAYER M1 ;
      RECT 1165 129695 1415 133225 ;
    LAYER M1 ;
      RECT 1165 133475 1415 134485 ;
    LAYER M1 ;
      RECT 1165 135575 1415 139105 ;
    LAYER M1 ;
      RECT 1165 139355 1415 140365 ;
    LAYER M1 ;
      RECT 1165 141455 1415 144985 ;
    LAYER M1 ;
      RECT 1165 145235 1415 146245 ;
    LAYER M1 ;
      RECT 1165 147335 1415 150865 ;
    LAYER M1 ;
      RECT 1165 151115 1415 152125 ;
    LAYER M1 ;
      RECT 1165 153215 1415 156745 ;
    LAYER M1 ;
      RECT 1165 156995 1415 158005 ;
    LAYER M1 ;
      RECT 1165 159095 1415 162625 ;
    LAYER M1 ;
      RECT 1165 162875 1415 163885 ;
    LAYER M1 ;
      RECT 1165 164975 1415 168505 ;
    LAYER M1 ;
      RECT 1165 168755 1415 169765 ;
    LAYER M1 ;
      RECT 1165 170855 1415 174385 ;
    LAYER M1 ;
      RECT 1165 174635 1415 175645 ;
    LAYER M1 ;
      RECT 1165 176735 1415 180265 ;
    LAYER M1 ;
      RECT 1165 180515 1415 181525 ;
    LAYER M1 ;
      RECT 1165 182615 1415 186145 ;
    LAYER M1 ;
      RECT 1165 186395 1415 187405 ;
    LAYER M1 ;
      RECT 1165 188495 1415 192025 ;
    LAYER M1 ;
      RECT 1165 192275 1415 193285 ;
    LAYER M1 ;
      RECT 1165 194375 1415 197905 ;
    LAYER M1 ;
      RECT 1165 198155 1415 199165 ;
    LAYER M1 ;
      RECT 1165 200255 1415 203785 ;
    LAYER M1 ;
      RECT 1165 204035 1415 205045 ;
    LAYER M1 ;
      RECT 1165 206135 1415 209665 ;
    LAYER M1 ;
      RECT 1165 209915 1415 210925 ;
    LAYER M1 ;
      RECT 1165 212015 1415 215545 ;
    LAYER M1 ;
      RECT 1165 215795 1415 216805 ;
    LAYER M1 ;
      RECT 1165 217895 1415 221425 ;
    LAYER M1 ;
      RECT 1165 221675 1415 222685 ;
    LAYER M1 ;
      RECT 1165 223775 1415 227305 ;
    LAYER M1 ;
      RECT 1165 227555 1415 228565 ;
    LAYER M1 ;
      RECT 1165 229655 1415 233185 ;
    LAYER M1 ;
      RECT 1165 233435 1415 234445 ;
    LAYER M1 ;
      RECT 1165 235535 1415 236545 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 735 59135 985 62665 ;
    LAYER M1 ;
      RECT 735 65015 985 68545 ;
    LAYER M1 ;
      RECT 735 70895 985 74425 ;
    LAYER M1 ;
      RECT 735 76775 985 80305 ;
    LAYER M1 ;
      RECT 735 82655 985 86185 ;
    LAYER M1 ;
      RECT 735 88535 985 92065 ;
    LAYER M1 ;
      RECT 735 94415 985 97945 ;
    LAYER M1 ;
      RECT 735 100295 985 103825 ;
    LAYER M1 ;
      RECT 735 106175 985 109705 ;
    LAYER M1 ;
      RECT 735 112055 985 115585 ;
    LAYER M1 ;
      RECT 735 117935 985 121465 ;
    LAYER M1 ;
      RECT 735 123815 985 127345 ;
    LAYER M1 ;
      RECT 735 129695 985 133225 ;
    LAYER M1 ;
      RECT 735 135575 985 139105 ;
    LAYER M1 ;
      RECT 735 141455 985 144985 ;
    LAYER M1 ;
      RECT 735 147335 985 150865 ;
    LAYER M1 ;
      RECT 735 153215 985 156745 ;
    LAYER M1 ;
      RECT 735 159095 985 162625 ;
    LAYER M1 ;
      RECT 735 164975 985 168505 ;
    LAYER M1 ;
      RECT 735 170855 985 174385 ;
    LAYER M1 ;
      RECT 735 176735 985 180265 ;
    LAYER M1 ;
      RECT 735 182615 985 186145 ;
    LAYER M1 ;
      RECT 735 188495 985 192025 ;
    LAYER M1 ;
      RECT 735 194375 985 197905 ;
    LAYER M1 ;
      RECT 735 200255 985 203785 ;
    LAYER M1 ;
      RECT 735 206135 985 209665 ;
    LAYER M1 ;
      RECT 735 212015 985 215545 ;
    LAYER M1 ;
      RECT 735 217895 985 221425 ;
    LAYER M1 ;
      RECT 735 223775 985 227305 ;
    LAYER M1 ;
      RECT 735 229655 985 233185 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M1 ;
      RECT 1595 59135 1845 62665 ;
    LAYER M1 ;
      RECT 1595 65015 1845 68545 ;
    LAYER M1 ;
      RECT 1595 70895 1845 74425 ;
    LAYER M1 ;
      RECT 1595 76775 1845 80305 ;
    LAYER M1 ;
      RECT 1595 82655 1845 86185 ;
    LAYER M1 ;
      RECT 1595 88535 1845 92065 ;
    LAYER M1 ;
      RECT 1595 94415 1845 97945 ;
    LAYER M1 ;
      RECT 1595 100295 1845 103825 ;
    LAYER M1 ;
      RECT 1595 106175 1845 109705 ;
    LAYER M1 ;
      RECT 1595 112055 1845 115585 ;
    LAYER M1 ;
      RECT 1595 117935 1845 121465 ;
    LAYER M1 ;
      RECT 1595 123815 1845 127345 ;
    LAYER M1 ;
      RECT 1595 129695 1845 133225 ;
    LAYER M1 ;
      RECT 1595 135575 1845 139105 ;
    LAYER M1 ;
      RECT 1595 141455 1845 144985 ;
    LAYER M1 ;
      RECT 1595 147335 1845 150865 ;
    LAYER M1 ;
      RECT 1595 153215 1845 156745 ;
    LAYER M1 ;
      RECT 1595 159095 1845 162625 ;
    LAYER M1 ;
      RECT 1595 164975 1845 168505 ;
    LAYER M1 ;
      RECT 1595 170855 1845 174385 ;
    LAYER M1 ;
      RECT 1595 176735 1845 180265 ;
    LAYER M1 ;
      RECT 1595 182615 1845 186145 ;
    LAYER M1 ;
      RECT 1595 188495 1845 192025 ;
    LAYER M1 ;
      RECT 1595 194375 1845 197905 ;
    LAYER M1 ;
      RECT 1595 200255 1845 203785 ;
    LAYER M1 ;
      RECT 1595 206135 1845 209665 ;
    LAYER M1 ;
      RECT 1595 212015 1845 215545 ;
    LAYER M1 ;
      RECT 1595 217895 1845 221425 ;
    LAYER M1 ;
      RECT 1595 223775 1845 227305 ;
    LAYER M1 ;
      RECT 1595 229655 1845 233185 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 33265 ;
    LAYER M1 ;
      RECT 2025 33515 2275 34525 ;
    LAYER M1 ;
      RECT 2025 35615 2275 39145 ;
    LAYER M1 ;
      RECT 2025 39395 2275 40405 ;
    LAYER M1 ;
      RECT 2025 41495 2275 45025 ;
    LAYER M1 ;
      RECT 2025 45275 2275 46285 ;
    LAYER M1 ;
      RECT 2025 47375 2275 50905 ;
    LAYER M1 ;
      RECT 2025 51155 2275 52165 ;
    LAYER M1 ;
      RECT 2025 53255 2275 56785 ;
    LAYER M1 ;
      RECT 2025 57035 2275 58045 ;
    LAYER M1 ;
      RECT 2025 59135 2275 62665 ;
    LAYER M1 ;
      RECT 2025 62915 2275 63925 ;
    LAYER M1 ;
      RECT 2025 65015 2275 68545 ;
    LAYER M1 ;
      RECT 2025 68795 2275 69805 ;
    LAYER M1 ;
      RECT 2025 70895 2275 74425 ;
    LAYER M1 ;
      RECT 2025 74675 2275 75685 ;
    LAYER M1 ;
      RECT 2025 76775 2275 80305 ;
    LAYER M1 ;
      RECT 2025 80555 2275 81565 ;
    LAYER M1 ;
      RECT 2025 82655 2275 86185 ;
    LAYER M1 ;
      RECT 2025 86435 2275 87445 ;
    LAYER M1 ;
      RECT 2025 88535 2275 92065 ;
    LAYER M1 ;
      RECT 2025 92315 2275 93325 ;
    LAYER M1 ;
      RECT 2025 94415 2275 97945 ;
    LAYER M1 ;
      RECT 2025 98195 2275 99205 ;
    LAYER M1 ;
      RECT 2025 100295 2275 103825 ;
    LAYER M1 ;
      RECT 2025 104075 2275 105085 ;
    LAYER M1 ;
      RECT 2025 106175 2275 109705 ;
    LAYER M1 ;
      RECT 2025 109955 2275 110965 ;
    LAYER M1 ;
      RECT 2025 112055 2275 115585 ;
    LAYER M1 ;
      RECT 2025 115835 2275 116845 ;
    LAYER M1 ;
      RECT 2025 117935 2275 121465 ;
    LAYER M1 ;
      RECT 2025 121715 2275 122725 ;
    LAYER M1 ;
      RECT 2025 123815 2275 127345 ;
    LAYER M1 ;
      RECT 2025 127595 2275 128605 ;
    LAYER M1 ;
      RECT 2025 129695 2275 133225 ;
    LAYER M1 ;
      RECT 2025 133475 2275 134485 ;
    LAYER M1 ;
      RECT 2025 135575 2275 139105 ;
    LAYER M1 ;
      RECT 2025 139355 2275 140365 ;
    LAYER M1 ;
      RECT 2025 141455 2275 144985 ;
    LAYER M1 ;
      RECT 2025 145235 2275 146245 ;
    LAYER M1 ;
      RECT 2025 147335 2275 150865 ;
    LAYER M1 ;
      RECT 2025 151115 2275 152125 ;
    LAYER M1 ;
      RECT 2025 153215 2275 156745 ;
    LAYER M1 ;
      RECT 2025 156995 2275 158005 ;
    LAYER M1 ;
      RECT 2025 159095 2275 162625 ;
    LAYER M1 ;
      RECT 2025 162875 2275 163885 ;
    LAYER M1 ;
      RECT 2025 164975 2275 168505 ;
    LAYER M1 ;
      RECT 2025 168755 2275 169765 ;
    LAYER M1 ;
      RECT 2025 170855 2275 174385 ;
    LAYER M1 ;
      RECT 2025 174635 2275 175645 ;
    LAYER M1 ;
      RECT 2025 176735 2275 180265 ;
    LAYER M1 ;
      RECT 2025 180515 2275 181525 ;
    LAYER M1 ;
      RECT 2025 182615 2275 186145 ;
    LAYER M1 ;
      RECT 2025 186395 2275 187405 ;
    LAYER M1 ;
      RECT 2025 188495 2275 192025 ;
    LAYER M1 ;
      RECT 2025 192275 2275 193285 ;
    LAYER M1 ;
      RECT 2025 194375 2275 197905 ;
    LAYER M1 ;
      RECT 2025 198155 2275 199165 ;
    LAYER M1 ;
      RECT 2025 200255 2275 203785 ;
    LAYER M1 ;
      RECT 2025 204035 2275 205045 ;
    LAYER M1 ;
      RECT 2025 206135 2275 209665 ;
    LAYER M1 ;
      RECT 2025 209915 2275 210925 ;
    LAYER M1 ;
      RECT 2025 212015 2275 215545 ;
    LAYER M1 ;
      RECT 2025 215795 2275 216805 ;
    LAYER M1 ;
      RECT 2025 217895 2275 221425 ;
    LAYER M1 ;
      RECT 2025 221675 2275 222685 ;
    LAYER M1 ;
      RECT 2025 223775 2275 227305 ;
    LAYER M1 ;
      RECT 2025 227555 2275 228565 ;
    LAYER M1 ;
      RECT 2025 229655 2275 233185 ;
    LAYER M1 ;
      RECT 2025 233435 2275 234445 ;
    LAYER M1 ;
      RECT 2025 235535 2275 236545 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2455 35615 2705 39145 ;
    LAYER M1 ;
      RECT 2455 41495 2705 45025 ;
    LAYER M1 ;
      RECT 2455 47375 2705 50905 ;
    LAYER M1 ;
      RECT 2455 53255 2705 56785 ;
    LAYER M1 ;
      RECT 2455 59135 2705 62665 ;
    LAYER M1 ;
      RECT 2455 65015 2705 68545 ;
    LAYER M1 ;
      RECT 2455 70895 2705 74425 ;
    LAYER M1 ;
      RECT 2455 76775 2705 80305 ;
    LAYER M1 ;
      RECT 2455 82655 2705 86185 ;
    LAYER M1 ;
      RECT 2455 88535 2705 92065 ;
    LAYER M1 ;
      RECT 2455 94415 2705 97945 ;
    LAYER M1 ;
      RECT 2455 100295 2705 103825 ;
    LAYER M1 ;
      RECT 2455 106175 2705 109705 ;
    LAYER M1 ;
      RECT 2455 112055 2705 115585 ;
    LAYER M1 ;
      RECT 2455 117935 2705 121465 ;
    LAYER M1 ;
      RECT 2455 123815 2705 127345 ;
    LAYER M1 ;
      RECT 2455 129695 2705 133225 ;
    LAYER M1 ;
      RECT 2455 135575 2705 139105 ;
    LAYER M1 ;
      RECT 2455 141455 2705 144985 ;
    LAYER M1 ;
      RECT 2455 147335 2705 150865 ;
    LAYER M1 ;
      RECT 2455 153215 2705 156745 ;
    LAYER M1 ;
      RECT 2455 159095 2705 162625 ;
    LAYER M1 ;
      RECT 2455 164975 2705 168505 ;
    LAYER M1 ;
      RECT 2455 170855 2705 174385 ;
    LAYER M1 ;
      RECT 2455 176735 2705 180265 ;
    LAYER M1 ;
      RECT 2455 182615 2705 186145 ;
    LAYER M1 ;
      RECT 2455 188495 2705 192025 ;
    LAYER M1 ;
      RECT 2455 194375 2705 197905 ;
    LAYER M1 ;
      RECT 2455 200255 2705 203785 ;
    LAYER M1 ;
      RECT 2455 206135 2705 209665 ;
    LAYER M1 ;
      RECT 2455 212015 2705 215545 ;
    LAYER M1 ;
      RECT 2455 217895 2705 221425 ;
    LAYER M1 ;
      RECT 2455 223775 2705 227305 ;
    LAYER M1 ;
      RECT 2455 229655 2705 233185 ;
    LAYER M2 ;
      RECT 1120 4480 2320 4760 ;
    LAYER M2 ;
      RECT 1120 280 2320 560 ;
    LAYER M2 ;
      RECT 690 700 2750 980 ;
    LAYER M2 ;
      RECT 1120 10360 2320 10640 ;
    LAYER M2 ;
      RECT 1120 6160 2320 6440 ;
    LAYER M2 ;
      RECT 690 6580 2750 6860 ;
    LAYER M2 ;
      RECT 1120 16240 2320 16520 ;
    LAYER M2 ;
      RECT 1120 12040 2320 12320 ;
    LAYER M2 ;
      RECT 690 12460 2750 12740 ;
    LAYER M2 ;
      RECT 1120 22120 2320 22400 ;
    LAYER M2 ;
      RECT 1120 17920 2320 18200 ;
    LAYER M2 ;
      RECT 690 18340 2750 18620 ;
    LAYER M2 ;
      RECT 1120 28000 2320 28280 ;
    LAYER M2 ;
      RECT 1120 23800 2320 24080 ;
    LAYER M2 ;
      RECT 690 24220 2750 24500 ;
    LAYER M2 ;
      RECT 1120 33880 2320 34160 ;
    LAYER M2 ;
      RECT 1120 29680 2320 29960 ;
    LAYER M2 ;
      RECT 690 30100 2750 30380 ;
    LAYER M2 ;
      RECT 1120 39760 2320 40040 ;
    LAYER M2 ;
      RECT 1120 35560 2320 35840 ;
    LAYER M2 ;
      RECT 690 35980 2750 36260 ;
    LAYER M2 ;
      RECT 1120 45640 2320 45920 ;
    LAYER M2 ;
      RECT 1120 41440 2320 41720 ;
    LAYER M2 ;
      RECT 690 41860 2750 42140 ;
    LAYER M2 ;
      RECT 1120 51520 2320 51800 ;
    LAYER M2 ;
      RECT 1120 47320 2320 47600 ;
    LAYER M2 ;
      RECT 690 47740 2750 48020 ;
    LAYER M2 ;
      RECT 1120 57400 2320 57680 ;
    LAYER M2 ;
      RECT 1120 53200 2320 53480 ;
    LAYER M2 ;
      RECT 690 53620 2750 53900 ;
    LAYER M2 ;
      RECT 1120 63280 2320 63560 ;
    LAYER M2 ;
      RECT 1120 59080 2320 59360 ;
    LAYER M2 ;
      RECT 690 59500 2750 59780 ;
    LAYER M2 ;
      RECT 1120 69160 2320 69440 ;
    LAYER M2 ;
      RECT 1120 64960 2320 65240 ;
    LAYER M2 ;
      RECT 690 65380 2750 65660 ;
    LAYER M2 ;
      RECT 1120 75040 2320 75320 ;
    LAYER M2 ;
      RECT 1120 70840 2320 71120 ;
    LAYER M2 ;
      RECT 690 71260 2750 71540 ;
    LAYER M2 ;
      RECT 1120 80920 2320 81200 ;
    LAYER M2 ;
      RECT 1120 76720 2320 77000 ;
    LAYER M2 ;
      RECT 690 77140 2750 77420 ;
    LAYER M2 ;
      RECT 1120 86800 2320 87080 ;
    LAYER M2 ;
      RECT 1120 82600 2320 82880 ;
    LAYER M2 ;
      RECT 690 83020 2750 83300 ;
    LAYER M2 ;
      RECT 1120 92680 2320 92960 ;
    LAYER M2 ;
      RECT 1120 88480 2320 88760 ;
    LAYER M2 ;
      RECT 690 88900 2750 89180 ;
    LAYER M2 ;
      RECT 1120 98560 2320 98840 ;
    LAYER M2 ;
      RECT 1120 94360 2320 94640 ;
    LAYER M2 ;
      RECT 690 94780 2750 95060 ;
    LAYER M2 ;
      RECT 1120 104440 2320 104720 ;
    LAYER M2 ;
      RECT 1120 100240 2320 100520 ;
    LAYER M2 ;
      RECT 690 100660 2750 100940 ;
    LAYER M2 ;
      RECT 1120 110320 2320 110600 ;
    LAYER M2 ;
      RECT 1120 106120 2320 106400 ;
    LAYER M2 ;
      RECT 690 106540 2750 106820 ;
    LAYER M2 ;
      RECT 1120 116200 2320 116480 ;
    LAYER M2 ;
      RECT 1120 112000 2320 112280 ;
    LAYER M2 ;
      RECT 690 112420 2750 112700 ;
    LAYER M2 ;
      RECT 1120 122080 2320 122360 ;
    LAYER M2 ;
      RECT 1120 117880 2320 118160 ;
    LAYER M2 ;
      RECT 690 118300 2750 118580 ;
    LAYER M2 ;
      RECT 1120 127960 2320 128240 ;
    LAYER M2 ;
      RECT 1120 123760 2320 124040 ;
    LAYER M2 ;
      RECT 690 124180 2750 124460 ;
    LAYER M2 ;
      RECT 1120 133840 2320 134120 ;
    LAYER M2 ;
      RECT 1120 129640 2320 129920 ;
    LAYER M2 ;
      RECT 690 130060 2750 130340 ;
    LAYER M2 ;
      RECT 1120 139720 2320 140000 ;
    LAYER M2 ;
      RECT 1120 135520 2320 135800 ;
    LAYER M2 ;
      RECT 690 135940 2750 136220 ;
    LAYER M2 ;
      RECT 1120 145600 2320 145880 ;
    LAYER M2 ;
      RECT 1120 141400 2320 141680 ;
    LAYER M2 ;
      RECT 690 141820 2750 142100 ;
    LAYER M2 ;
      RECT 1120 151480 2320 151760 ;
    LAYER M2 ;
      RECT 1120 147280 2320 147560 ;
    LAYER M2 ;
      RECT 690 147700 2750 147980 ;
    LAYER M2 ;
      RECT 1120 157360 2320 157640 ;
    LAYER M2 ;
      RECT 1120 153160 2320 153440 ;
    LAYER M2 ;
      RECT 690 153580 2750 153860 ;
    LAYER M2 ;
      RECT 1120 163240 2320 163520 ;
    LAYER M2 ;
      RECT 1120 159040 2320 159320 ;
    LAYER M2 ;
      RECT 690 159460 2750 159740 ;
    LAYER M2 ;
      RECT 1120 169120 2320 169400 ;
    LAYER M2 ;
      RECT 1120 164920 2320 165200 ;
    LAYER M2 ;
      RECT 690 165340 2750 165620 ;
    LAYER M2 ;
      RECT 1120 175000 2320 175280 ;
    LAYER M2 ;
      RECT 1120 170800 2320 171080 ;
    LAYER M2 ;
      RECT 690 171220 2750 171500 ;
    LAYER M2 ;
      RECT 1120 180880 2320 181160 ;
    LAYER M2 ;
      RECT 1120 176680 2320 176960 ;
    LAYER M2 ;
      RECT 690 177100 2750 177380 ;
    LAYER M2 ;
      RECT 1120 186760 2320 187040 ;
    LAYER M2 ;
      RECT 1120 182560 2320 182840 ;
    LAYER M2 ;
      RECT 690 182980 2750 183260 ;
    LAYER M2 ;
      RECT 1120 192640 2320 192920 ;
    LAYER M2 ;
      RECT 1120 188440 2320 188720 ;
    LAYER M2 ;
      RECT 690 188860 2750 189140 ;
    LAYER M2 ;
      RECT 1120 198520 2320 198800 ;
    LAYER M2 ;
      RECT 1120 194320 2320 194600 ;
    LAYER M2 ;
      RECT 690 194740 2750 195020 ;
    LAYER M2 ;
      RECT 1120 204400 2320 204680 ;
    LAYER M2 ;
      RECT 1120 200200 2320 200480 ;
    LAYER M2 ;
      RECT 690 200620 2750 200900 ;
    LAYER M2 ;
      RECT 1120 210280 2320 210560 ;
    LAYER M2 ;
      RECT 1120 206080 2320 206360 ;
    LAYER M2 ;
      RECT 690 206500 2750 206780 ;
    LAYER M2 ;
      RECT 1120 216160 2320 216440 ;
    LAYER M2 ;
      RECT 1120 211960 2320 212240 ;
    LAYER M2 ;
      RECT 690 212380 2750 212660 ;
    LAYER M2 ;
      RECT 1120 222040 2320 222320 ;
    LAYER M2 ;
      RECT 1120 217840 2320 218120 ;
    LAYER M2 ;
      RECT 690 218260 2750 218540 ;
    LAYER M2 ;
      RECT 1120 227920 2320 228200 ;
    LAYER M2 ;
      RECT 1120 223720 2320 224000 ;
    LAYER M2 ;
      RECT 690 224140 2750 224420 ;
    LAYER M2 ;
      RECT 1120 233800 2320 234080 ;
    LAYER M2 ;
      RECT 1120 229600 2320 229880 ;
    LAYER M2 ;
      RECT 1120 235900 2320 236180 ;
    LAYER M2 ;
      RECT 690 230020 2750 230300 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53255 1375 53425 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59135 1375 59305 ;
    LAYER V1 ;
      RECT 1205 63335 1375 63505 ;
    LAYER V1 ;
      RECT 1205 65015 1375 65185 ;
    LAYER V1 ;
      RECT 1205 69215 1375 69385 ;
    LAYER V1 ;
      RECT 1205 70895 1375 71065 ;
    LAYER V1 ;
      RECT 1205 75095 1375 75265 ;
    LAYER V1 ;
      RECT 1205 76775 1375 76945 ;
    LAYER V1 ;
      RECT 1205 80975 1375 81145 ;
    LAYER V1 ;
      RECT 1205 82655 1375 82825 ;
    LAYER V1 ;
      RECT 1205 86855 1375 87025 ;
    LAYER V1 ;
      RECT 1205 88535 1375 88705 ;
    LAYER V1 ;
      RECT 1205 92735 1375 92905 ;
    LAYER V1 ;
      RECT 1205 94415 1375 94585 ;
    LAYER V1 ;
      RECT 1205 98615 1375 98785 ;
    LAYER V1 ;
      RECT 1205 100295 1375 100465 ;
    LAYER V1 ;
      RECT 1205 104495 1375 104665 ;
    LAYER V1 ;
      RECT 1205 106175 1375 106345 ;
    LAYER V1 ;
      RECT 1205 110375 1375 110545 ;
    LAYER V1 ;
      RECT 1205 112055 1375 112225 ;
    LAYER V1 ;
      RECT 1205 116255 1375 116425 ;
    LAYER V1 ;
      RECT 1205 117935 1375 118105 ;
    LAYER V1 ;
      RECT 1205 122135 1375 122305 ;
    LAYER V1 ;
      RECT 1205 123815 1375 123985 ;
    LAYER V1 ;
      RECT 1205 128015 1375 128185 ;
    LAYER V1 ;
      RECT 1205 129695 1375 129865 ;
    LAYER V1 ;
      RECT 1205 133895 1375 134065 ;
    LAYER V1 ;
      RECT 1205 135575 1375 135745 ;
    LAYER V1 ;
      RECT 1205 139775 1375 139945 ;
    LAYER V1 ;
      RECT 1205 141455 1375 141625 ;
    LAYER V1 ;
      RECT 1205 145655 1375 145825 ;
    LAYER V1 ;
      RECT 1205 147335 1375 147505 ;
    LAYER V1 ;
      RECT 1205 151535 1375 151705 ;
    LAYER V1 ;
      RECT 1205 153215 1375 153385 ;
    LAYER V1 ;
      RECT 1205 157415 1375 157585 ;
    LAYER V1 ;
      RECT 1205 159095 1375 159265 ;
    LAYER V1 ;
      RECT 1205 163295 1375 163465 ;
    LAYER V1 ;
      RECT 1205 164975 1375 165145 ;
    LAYER V1 ;
      RECT 1205 169175 1375 169345 ;
    LAYER V1 ;
      RECT 1205 170855 1375 171025 ;
    LAYER V1 ;
      RECT 1205 175055 1375 175225 ;
    LAYER V1 ;
      RECT 1205 176735 1375 176905 ;
    LAYER V1 ;
      RECT 1205 180935 1375 181105 ;
    LAYER V1 ;
      RECT 1205 182615 1375 182785 ;
    LAYER V1 ;
      RECT 1205 186815 1375 186985 ;
    LAYER V1 ;
      RECT 1205 188495 1375 188665 ;
    LAYER V1 ;
      RECT 1205 192695 1375 192865 ;
    LAYER V1 ;
      RECT 1205 194375 1375 194545 ;
    LAYER V1 ;
      RECT 1205 198575 1375 198745 ;
    LAYER V1 ;
      RECT 1205 200255 1375 200425 ;
    LAYER V1 ;
      RECT 1205 204455 1375 204625 ;
    LAYER V1 ;
      RECT 1205 206135 1375 206305 ;
    LAYER V1 ;
      RECT 1205 210335 1375 210505 ;
    LAYER V1 ;
      RECT 1205 212015 1375 212185 ;
    LAYER V1 ;
      RECT 1205 216215 1375 216385 ;
    LAYER V1 ;
      RECT 1205 217895 1375 218065 ;
    LAYER V1 ;
      RECT 1205 222095 1375 222265 ;
    LAYER V1 ;
      RECT 1205 223775 1375 223945 ;
    LAYER V1 ;
      RECT 1205 227975 1375 228145 ;
    LAYER V1 ;
      RECT 1205 229655 1375 229825 ;
    LAYER V1 ;
      RECT 1205 233855 1375 234025 ;
    LAYER V1 ;
      RECT 1205 235955 1375 236125 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 29735 2235 29905 ;
    LAYER V1 ;
      RECT 2065 33935 2235 34105 ;
    LAYER V1 ;
      RECT 2065 35615 2235 35785 ;
    LAYER V1 ;
      RECT 2065 39815 2235 39985 ;
    LAYER V1 ;
      RECT 2065 41495 2235 41665 ;
    LAYER V1 ;
      RECT 2065 45695 2235 45865 ;
    LAYER V1 ;
      RECT 2065 47375 2235 47545 ;
    LAYER V1 ;
      RECT 2065 51575 2235 51745 ;
    LAYER V1 ;
      RECT 2065 53255 2235 53425 ;
    LAYER V1 ;
      RECT 2065 57455 2235 57625 ;
    LAYER V1 ;
      RECT 2065 59135 2235 59305 ;
    LAYER V1 ;
      RECT 2065 63335 2235 63505 ;
    LAYER V1 ;
      RECT 2065 65015 2235 65185 ;
    LAYER V1 ;
      RECT 2065 69215 2235 69385 ;
    LAYER V1 ;
      RECT 2065 70895 2235 71065 ;
    LAYER V1 ;
      RECT 2065 75095 2235 75265 ;
    LAYER V1 ;
      RECT 2065 76775 2235 76945 ;
    LAYER V1 ;
      RECT 2065 80975 2235 81145 ;
    LAYER V1 ;
      RECT 2065 82655 2235 82825 ;
    LAYER V1 ;
      RECT 2065 86855 2235 87025 ;
    LAYER V1 ;
      RECT 2065 88535 2235 88705 ;
    LAYER V1 ;
      RECT 2065 92735 2235 92905 ;
    LAYER V1 ;
      RECT 2065 94415 2235 94585 ;
    LAYER V1 ;
      RECT 2065 98615 2235 98785 ;
    LAYER V1 ;
      RECT 2065 100295 2235 100465 ;
    LAYER V1 ;
      RECT 2065 104495 2235 104665 ;
    LAYER V1 ;
      RECT 2065 106175 2235 106345 ;
    LAYER V1 ;
      RECT 2065 110375 2235 110545 ;
    LAYER V1 ;
      RECT 2065 112055 2235 112225 ;
    LAYER V1 ;
      RECT 2065 116255 2235 116425 ;
    LAYER V1 ;
      RECT 2065 117935 2235 118105 ;
    LAYER V1 ;
      RECT 2065 122135 2235 122305 ;
    LAYER V1 ;
      RECT 2065 123815 2235 123985 ;
    LAYER V1 ;
      RECT 2065 128015 2235 128185 ;
    LAYER V1 ;
      RECT 2065 129695 2235 129865 ;
    LAYER V1 ;
      RECT 2065 133895 2235 134065 ;
    LAYER V1 ;
      RECT 2065 135575 2235 135745 ;
    LAYER V1 ;
      RECT 2065 139775 2235 139945 ;
    LAYER V1 ;
      RECT 2065 141455 2235 141625 ;
    LAYER V1 ;
      RECT 2065 145655 2235 145825 ;
    LAYER V1 ;
      RECT 2065 147335 2235 147505 ;
    LAYER V1 ;
      RECT 2065 151535 2235 151705 ;
    LAYER V1 ;
      RECT 2065 153215 2235 153385 ;
    LAYER V1 ;
      RECT 2065 157415 2235 157585 ;
    LAYER V1 ;
      RECT 2065 159095 2235 159265 ;
    LAYER V1 ;
      RECT 2065 163295 2235 163465 ;
    LAYER V1 ;
      RECT 2065 164975 2235 165145 ;
    LAYER V1 ;
      RECT 2065 169175 2235 169345 ;
    LAYER V1 ;
      RECT 2065 170855 2235 171025 ;
    LAYER V1 ;
      RECT 2065 175055 2235 175225 ;
    LAYER V1 ;
      RECT 2065 176735 2235 176905 ;
    LAYER V1 ;
      RECT 2065 180935 2235 181105 ;
    LAYER V1 ;
      RECT 2065 182615 2235 182785 ;
    LAYER V1 ;
      RECT 2065 186815 2235 186985 ;
    LAYER V1 ;
      RECT 2065 188495 2235 188665 ;
    LAYER V1 ;
      RECT 2065 192695 2235 192865 ;
    LAYER V1 ;
      RECT 2065 194375 2235 194545 ;
    LAYER V1 ;
      RECT 2065 198575 2235 198745 ;
    LAYER V1 ;
      RECT 2065 200255 2235 200425 ;
    LAYER V1 ;
      RECT 2065 204455 2235 204625 ;
    LAYER V1 ;
      RECT 2065 206135 2235 206305 ;
    LAYER V1 ;
      RECT 2065 210335 2235 210505 ;
    LAYER V1 ;
      RECT 2065 212015 2235 212185 ;
    LAYER V1 ;
      RECT 2065 216215 2235 216385 ;
    LAYER V1 ;
      RECT 2065 217895 2235 218065 ;
    LAYER V1 ;
      RECT 2065 222095 2235 222265 ;
    LAYER V1 ;
      RECT 2065 223775 2235 223945 ;
    LAYER V1 ;
      RECT 2065 227975 2235 228145 ;
    LAYER V1 ;
      RECT 2065 229655 2235 229825 ;
    LAYER V1 ;
      RECT 2065 233855 2235 234025 ;
    LAYER V1 ;
      RECT 2065 235955 2235 236125 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 775 53675 945 53845 ;
    LAYER V1 ;
      RECT 775 59555 945 59725 ;
    LAYER V1 ;
      RECT 775 65435 945 65605 ;
    LAYER V1 ;
      RECT 775 71315 945 71485 ;
    LAYER V1 ;
      RECT 775 77195 945 77365 ;
    LAYER V1 ;
      RECT 775 83075 945 83245 ;
    LAYER V1 ;
      RECT 775 88955 945 89125 ;
    LAYER V1 ;
      RECT 775 94835 945 95005 ;
    LAYER V1 ;
      RECT 775 100715 945 100885 ;
    LAYER V1 ;
      RECT 775 106595 945 106765 ;
    LAYER V1 ;
      RECT 775 112475 945 112645 ;
    LAYER V1 ;
      RECT 775 118355 945 118525 ;
    LAYER V1 ;
      RECT 775 124235 945 124405 ;
    LAYER V1 ;
      RECT 775 130115 945 130285 ;
    LAYER V1 ;
      RECT 775 135995 945 136165 ;
    LAYER V1 ;
      RECT 775 141875 945 142045 ;
    LAYER V1 ;
      RECT 775 147755 945 147925 ;
    LAYER V1 ;
      RECT 775 153635 945 153805 ;
    LAYER V1 ;
      RECT 775 159515 945 159685 ;
    LAYER V1 ;
      RECT 775 165395 945 165565 ;
    LAYER V1 ;
      RECT 775 171275 945 171445 ;
    LAYER V1 ;
      RECT 775 177155 945 177325 ;
    LAYER V1 ;
      RECT 775 183035 945 183205 ;
    LAYER V1 ;
      RECT 775 188915 945 189085 ;
    LAYER V1 ;
      RECT 775 194795 945 194965 ;
    LAYER V1 ;
      RECT 775 200675 945 200845 ;
    LAYER V1 ;
      RECT 775 206555 945 206725 ;
    LAYER V1 ;
      RECT 775 212435 945 212605 ;
    LAYER V1 ;
      RECT 775 218315 945 218485 ;
    LAYER V1 ;
      RECT 775 224195 945 224365 ;
    LAYER V1 ;
      RECT 775 230075 945 230245 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 1635 53675 1805 53845 ;
    LAYER V1 ;
      RECT 1635 59555 1805 59725 ;
    LAYER V1 ;
      RECT 1635 65435 1805 65605 ;
    LAYER V1 ;
      RECT 1635 71315 1805 71485 ;
    LAYER V1 ;
      RECT 1635 77195 1805 77365 ;
    LAYER V1 ;
      RECT 1635 83075 1805 83245 ;
    LAYER V1 ;
      RECT 1635 88955 1805 89125 ;
    LAYER V1 ;
      RECT 1635 94835 1805 95005 ;
    LAYER V1 ;
      RECT 1635 100715 1805 100885 ;
    LAYER V1 ;
      RECT 1635 106595 1805 106765 ;
    LAYER V1 ;
      RECT 1635 112475 1805 112645 ;
    LAYER V1 ;
      RECT 1635 118355 1805 118525 ;
    LAYER V1 ;
      RECT 1635 124235 1805 124405 ;
    LAYER V1 ;
      RECT 1635 130115 1805 130285 ;
    LAYER V1 ;
      RECT 1635 135995 1805 136165 ;
    LAYER V1 ;
      RECT 1635 141875 1805 142045 ;
    LAYER V1 ;
      RECT 1635 147755 1805 147925 ;
    LAYER V1 ;
      RECT 1635 153635 1805 153805 ;
    LAYER V1 ;
      RECT 1635 159515 1805 159685 ;
    LAYER V1 ;
      RECT 1635 165395 1805 165565 ;
    LAYER V1 ;
      RECT 1635 171275 1805 171445 ;
    LAYER V1 ;
      RECT 1635 177155 1805 177325 ;
    LAYER V1 ;
      RECT 1635 183035 1805 183205 ;
    LAYER V1 ;
      RECT 1635 188915 1805 189085 ;
    LAYER V1 ;
      RECT 1635 194795 1805 194965 ;
    LAYER V1 ;
      RECT 1635 200675 1805 200845 ;
    LAYER V1 ;
      RECT 1635 206555 1805 206725 ;
    LAYER V1 ;
      RECT 1635 212435 1805 212605 ;
    LAYER V1 ;
      RECT 1635 218315 1805 218485 ;
    LAYER V1 ;
      RECT 1635 224195 1805 224365 ;
    LAYER V1 ;
      RECT 1635 230075 1805 230245 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 2495 30155 2665 30325 ;
    LAYER V1 ;
      RECT 2495 36035 2665 36205 ;
    LAYER V1 ;
      RECT 2495 41915 2665 42085 ;
    LAYER V1 ;
      RECT 2495 47795 2665 47965 ;
    LAYER V1 ;
      RECT 2495 53675 2665 53845 ;
    LAYER V1 ;
      RECT 2495 59555 2665 59725 ;
    LAYER V1 ;
      RECT 2495 65435 2665 65605 ;
    LAYER V1 ;
      RECT 2495 71315 2665 71485 ;
    LAYER V1 ;
      RECT 2495 77195 2665 77365 ;
    LAYER V1 ;
      RECT 2495 83075 2665 83245 ;
    LAYER V1 ;
      RECT 2495 88955 2665 89125 ;
    LAYER V1 ;
      RECT 2495 94835 2665 95005 ;
    LAYER V1 ;
      RECT 2495 100715 2665 100885 ;
    LAYER V1 ;
      RECT 2495 106595 2665 106765 ;
    LAYER V1 ;
      RECT 2495 112475 2665 112645 ;
    LAYER V1 ;
      RECT 2495 118355 2665 118525 ;
    LAYER V1 ;
      RECT 2495 124235 2665 124405 ;
    LAYER V1 ;
      RECT 2495 130115 2665 130285 ;
    LAYER V1 ;
      RECT 2495 135995 2665 136165 ;
    LAYER V1 ;
      RECT 2495 141875 2665 142045 ;
    LAYER V1 ;
      RECT 2495 147755 2665 147925 ;
    LAYER V1 ;
      RECT 2495 153635 2665 153805 ;
    LAYER V1 ;
      RECT 2495 159515 2665 159685 ;
    LAYER V1 ;
      RECT 2495 165395 2665 165565 ;
    LAYER V1 ;
      RECT 2495 171275 2665 171445 ;
    LAYER V1 ;
      RECT 2495 177155 2665 177325 ;
    LAYER V1 ;
      RECT 2495 183035 2665 183205 ;
    LAYER V1 ;
      RECT 2495 188915 2665 189085 ;
    LAYER V1 ;
      RECT 2495 194795 2665 194965 ;
    LAYER V1 ;
      RECT 2495 200675 2665 200845 ;
    LAYER V1 ;
      RECT 2495 206555 2665 206725 ;
    LAYER V1 ;
      RECT 2495 212435 2665 212605 ;
    LAYER V1 ;
      RECT 2495 218315 2665 218485 ;
    LAYER V1 ;
      RECT 2495 224195 2665 224365 ;
    LAYER V1 ;
      RECT 2495 230075 2665 230245 ;
    LAYER V2 ;
      RECT 1645 345 1795 495 ;
    LAYER V2 ;
      RECT 1645 4545 1795 4695 ;
    LAYER V2 ;
      RECT 1645 6225 1795 6375 ;
    LAYER V2 ;
      RECT 1645 10425 1795 10575 ;
    LAYER V2 ;
      RECT 1645 12105 1795 12255 ;
    LAYER V2 ;
      RECT 1645 16305 1795 16455 ;
    LAYER V2 ;
      RECT 1645 17985 1795 18135 ;
    LAYER V2 ;
      RECT 1645 22185 1795 22335 ;
    LAYER V2 ;
      RECT 1645 23865 1795 24015 ;
    LAYER V2 ;
      RECT 1645 28065 1795 28215 ;
    LAYER V2 ;
      RECT 1645 29745 1795 29895 ;
    LAYER V2 ;
      RECT 1645 33945 1795 34095 ;
    LAYER V2 ;
      RECT 1645 35625 1795 35775 ;
    LAYER V2 ;
      RECT 1645 39825 1795 39975 ;
    LAYER V2 ;
      RECT 1645 41505 1795 41655 ;
    LAYER V2 ;
      RECT 1645 45705 1795 45855 ;
    LAYER V2 ;
      RECT 1645 47385 1795 47535 ;
    LAYER V2 ;
      RECT 1645 51585 1795 51735 ;
    LAYER V2 ;
      RECT 1645 53265 1795 53415 ;
    LAYER V2 ;
      RECT 1645 57465 1795 57615 ;
    LAYER V2 ;
      RECT 1645 59145 1795 59295 ;
    LAYER V2 ;
      RECT 1645 63345 1795 63495 ;
    LAYER V2 ;
      RECT 1645 65025 1795 65175 ;
    LAYER V2 ;
      RECT 1645 69225 1795 69375 ;
    LAYER V2 ;
      RECT 1645 70905 1795 71055 ;
    LAYER V2 ;
      RECT 1645 75105 1795 75255 ;
    LAYER V2 ;
      RECT 1645 76785 1795 76935 ;
    LAYER V2 ;
      RECT 1645 80985 1795 81135 ;
    LAYER V2 ;
      RECT 1645 82665 1795 82815 ;
    LAYER V2 ;
      RECT 1645 86865 1795 87015 ;
    LAYER V2 ;
      RECT 1645 88545 1795 88695 ;
    LAYER V2 ;
      RECT 1645 92745 1795 92895 ;
    LAYER V2 ;
      RECT 1645 94425 1795 94575 ;
    LAYER V2 ;
      RECT 1645 98625 1795 98775 ;
    LAYER V2 ;
      RECT 1645 100305 1795 100455 ;
    LAYER V2 ;
      RECT 1645 104505 1795 104655 ;
    LAYER V2 ;
      RECT 1645 106185 1795 106335 ;
    LAYER V2 ;
      RECT 1645 110385 1795 110535 ;
    LAYER V2 ;
      RECT 1645 112065 1795 112215 ;
    LAYER V2 ;
      RECT 1645 116265 1795 116415 ;
    LAYER V2 ;
      RECT 1645 117945 1795 118095 ;
    LAYER V2 ;
      RECT 1645 122145 1795 122295 ;
    LAYER V2 ;
      RECT 1645 123825 1795 123975 ;
    LAYER V2 ;
      RECT 1645 128025 1795 128175 ;
    LAYER V2 ;
      RECT 1645 129705 1795 129855 ;
    LAYER V2 ;
      RECT 1645 133905 1795 134055 ;
    LAYER V2 ;
      RECT 1645 135585 1795 135735 ;
    LAYER V2 ;
      RECT 1645 139785 1795 139935 ;
    LAYER V2 ;
      RECT 1645 141465 1795 141615 ;
    LAYER V2 ;
      RECT 1645 145665 1795 145815 ;
    LAYER V2 ;
      RECT 1645 147345 1795 147495 ;
    LAYER V2 ;
      RECT 1645 151545 1795 151695 ;
    LAYER V2 ;
      RECT 1645 153225 1795 153375 ;
    LAYER V2 ;
      RECT 1645 157425 1795 157575 ;
    LAYER V2 ;
      RECT 1645 159105 1795 159255 ;
    LAYER V2 ;
      RECT 1645 163305 1795 163455 ;
    LAYER V2 ;
      RECT 1645 164985 1795 165135 ;
    LAYER V2 ;
      RECT 1645 169185 1795 169335 ;
    LAYER V2 ;
      RECT 1645 170865 1795 171015 ;
    LAYER V2 ;
      RECT 1645 175065 1795 175215 ;
    LAYER V2 ;
      RECT 1645 176745 1795 176895 ;
    LAYER V2 ;
      RECT 1645 180945 1795 181095 ;
    LAYER V2 ;
      RECT 1645 182625 1795 182775 ;
    LAYER V2 ;
      RECT 1645 186825 1795 186975 ;
    LAYER V2 ;
      RECT 1645 188505 1795 188655 ;
    LAYER V2 ;
      RECT 1645 192705 1795 192855 ;
    LAYER V2 ;
      RECT 1645 194385 1795 194535 ;
    LAYER V2 ;
      RECT 1645 198585 1795 198735 ;
    LAYER V2 ;
      RECT 1645 200265 1795 200415 ;
    LAYER V2 ;
      RECT 1645 204465 1795 204615 ;
    LAYER V2 ;
      RECT 1645 206145 1795 206295 ;
    LAYER V2 ;
      RECT 1645 210345 1795 210495 ;
    LAYER V2 ;
      RECT 1645 212025 1795 212175 ;
    LAYER V2 ;
      RECT 1645 216225 1795 216375 ;
    LAYER V2 ;
      RECT 1645 217905 1795 218055 ;
    LAYER V2 ;
      RECT 1645 222105 1795 222255 ;
    LAYER V2 ;
      RECT 1645 223785 1795 223935 ;
    LAYER V2 ;
      RECT 1645 227985 1795 228135 ;
    LAYER V2 ;
      RECT 1645 229665 1795 229815 ;
    LAYER V2 ;
      RECT 1645 233865 1795 234015 ;
    LAYER V2 ;
      RECT 2075 765 2225 915 ;
    LAYER V2 ;
      RECT 2075 6645 2225 6795 ;
    LAYER V2 ;
      RECT 2075 12525 2225 12675 ;
    LAYER V2 ;
      RECT 2075 18405 2225 18555 ;
    LAYER V2 ;
      RECT 2075 24285 2225 24435 ;
    LAYER V2 ;
      RECT 2075 30165 2225 30315 ;
    LAYER V2 ;
      RECT 2075 36045 2225 36195 ;
    LAYER V2 ;
      RECT 2075 41925 2225 42075 ;
    LAYER V2 ;
      RECT 2075 47805 2225 47955 ;
    LAYER V2 ;
      RECT 2075 53685 2225 53835 ;
    LAYER V2 ;
      RECT 2075 59565 2225 59715 ;
    LAYER V2 ;
      RECT 2075 65445 2225 65595 ;
    LAYER V2 ;
      RECT 2075 71325 2225 71475 ;
    LAYER V2 ;
      RECT 2075 77205 2225 77355 ;
    LAYER V2 ;
      RECT 2075 83085 2225 83235 ;
    LAYER V2 ;
      RECT 2075 88965 2225 89115 ;
    LAYER V2 ;
      RECT 2075 94845 2225 94995 ;
    LAYER V2 ;
      RECT 2075 100725 2225 100875 ;
    LAYER V2 ;
      RECT 2075 106605 2225 106755 ;
    LAYER V2 ;
      RECT 2075 112485 2225 112635 ;
    LAYER V2 ;
      RECT 2075 118365 2225 118515 ;
    LAYER V2 ;
      RECT 2075 124245 2225 124395 ;
    LAYER V2 ;
      RECT 2075 130125 2225 130275 ;
    LAYER V2 ;
      RECT 2075 136005 2225 136155 ;
    LAYER V2 ;
      RECT 2075 141885 2225 142035 ;
    LAYER V2 ;
      RECT 2075 147765 2225 147915 ;
    LAYER V2 ;
      RECT 2075 153645 2225 153795 ;
    LAYER V2 ;
      RECT 2075 159525 2225 159675 ;
    LAYER V2 ;
      RECT 2075 165405 2225 165555 ;
    LAYER V2 ;
      RECT 2075 171285 2225 171435 ;
    LAYER V2 ;
      RECT 2075 177165 2225 177315 ;
    LAYER V2 ;
      RECT 2075 183045 2225 183195 ;
    LAYER V2 ;
      RECT 2075 188925 2225 189075 ;
    LAYER V2 ;
      RECT 2075 194805 2225 194955 ;
    LAYER V2 ;
      RECT 2075 200685 2225 200835 ;
    LAYER V2 ;
      RECT 2075 206565 2225 206715 ;
    LAYER V2 ;
      RECT 2075 212445 2225 212595 ;
    LAYER V2 ;
      RECT 2075 218325 2225 218475 ;
    LAYER V2 ;
      RECT 2075 224205 2225 224355 ;
    LAYER V2 ;
      RECT 2075 230085 2225 230235 ;
    LAYER V2 ;
      RECT 2075 235965 2225 236115 ;
  END
END DCL_NMOS_S_42410075_X2_Y40
