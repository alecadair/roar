MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 53.91 BY 21.59 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 25.23 7.82 25.51 12.34 ;
      LAYER M2 ;
        RECT 26.92 12.04 28.12 12.32 ;
      LAYER M3 ;
        RECT 25.23 11.575 25.51 11.945 ;
      LAYER M2 ;
        RECT 25.37 11.62 27.09 11.9 ;
      LAYER M1 ;
        RECT 26.965 11.76 27.215 12.18 ;
      LAYER M2 ;
        RECT 26.93 12.04 27.25 12.32 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 12.33 6.98 12.61 13.18 ;
      LAYER M2 ;
        RECT 5.42 13.72 16.94 14 ;
      LAYER M3 ;
        RECT 12.33 13.02 12.61 13.86 ;
      LAYER M2 ;
        RECT 12.31 13.72 12.63 14 ;
    END
  END VOUT
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 24.34 2.8 25.54 3.08 ;
    END
  END VINN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 27.78 2.8 28.98 3.08 ;
    END
  END VINP
  OBS 
  LAYER M2 ;
        RECT 5.42 17.92 16.94 18.2 ;
  LAYER M3 ;
        RECT 42 13.7 42.28 18.22 ;
  LAYER M3 ;
        RECT 40.71 6.98 40.99 13.18 ;
  LAYER M2 ;
        RECT 16.77 17.92 18.49 18.2 ;
  LAYER M3 ;
        RECT 18.35 17.64 18.63 18.06 ;
  LAYER M2 ;
        RECT 18.49 17.5 42.14 17.78 ;
  LAYER M3 ;
        RECT 42 17.455 42.28 17.825 ;
  LAYER M3 ;
        RECT 42 13.675 42.28 14.045 ;
  LAYER M4 ;
        RECT 40.85 13.46 42.14 14.26 ;
  LAYER M3 ;
        RECT 40.71 13.02 40.99 13.86 ;
  LAYER M2 ;
        RECT 18.33 17.5 18.65 17.78 ;
  LAYER M3 ;
        RECT 18.35 17.48 18.63 17.8 ;
  LAYER M2 ;
        RECT 18.33 17.92 18.65 18.2 ;
  LAYER M3 ;
        RECT 18.35 17.9 18.63 18.22 ;
  LAYER M2 ;
        RECT 41.98 17.5 42.3 17.78 ;
  LAYER M3 ;
        RECT 42 17.48 42.28 17.8 ;
  LAYER M2 ;
        RECT 18.33 17.5 18.65 17.78 ;
  LAYER M3 ;
        RECT 18.35 17.48 18.63 17.8 ;
  LAYER M2 ;
        RECT 18.33 17.92 18.65 18.2 ;
  LAYER M3 ;
        RECT 18.35 17.9 18.63 18.22 ;
  LAYER M2 ;
        RECT 41.98 17.5 42.3 17.78 ;
  LAYER M3 ;
        RECT 42 17.48 42.28 17.8 ;
  LAYER M2 ;
        RECT 18.33 17.5 18.65 17.78 ;
  LAYER M3 ;
        RECT 18.35 17.48 18.63 17.8 ;
  LAYER M2 ;
        RECT 18.33 17.92 18.65 18.2 ;
  LAYER M3 ;
        RECT 18.35 17.9 18.63 18.22 ;
  LAYER M2 ;
        RECT 41.98 17.5 42.3 17.78 ;
  LAYER M3 ;
        RECT 42 17.48 42.28 17.8 ;
  LAYER M3 ;
        RECT 40.71 13.675 40.99 14.045 ;
  LAYER M4 ;
        RECT 40.685 13.46 41.015 14.26 ;
  LAYER M3 ;
        RECT 42 13.675 42.28 14.045 ;
  LAYER M4 ;
        RECT 41.975 13.46 42.305 14.26 ;
  LAYER M2 ;
        RECT 18.33 17.5 18.65 17.78 ;
  LAYER M3 ;
        RECT 18.35 17.48 18.63 17.8 ;
  LAYER M2 ;
        RECT 18.33 17.92 18.65 18.2 ;
  LAYER M3 ;
        RECT 18.35 17.9 18.63 18.22 ;
  LAYER M2 ;
        RECT 41.98 17.5 42.3 17.78 ;
  LAYER M3 ;
        RECT 42 17.48 42.28 17.8 ;
  LAYER M3 ;
        RECT 40.71 13.675 40.99 14.045 ;
  LAYER M4 ;
        RECT 40.685 13.46 41.015 14.26 ;
  LAYER M3 ;
        RECT 42 13.675 42.28 14.045 ;
  LAYER M4 ;
        RECT 41.975 13.46 42.305 14.26 ;
  LAYER M3 ;
        RECT 11.9 2.78 12.18 8.98 ;
  LAYER M2 ;
        RECT 24.34 7 25.54 7.28 ;
  LAYER M3 ;
        RECT 20.93 13.7 21.21 18.22 ;
  LAYER M3 ;
        RECT 11.9 7.375 12.18 7.745 ;
  LAYER M2 ;
        RECT 12.04 7.42 23.65 7.7 ;
  LAYER M1 ;
        RECT 23.525 7.14 23.775 7.56 ;
  LAYER M2 ;
        RECT 23.65 7 24.51 7.28 ;
  LAYER M2 ;
        RECT 20.91 7.42 21.23 7.7 ;
  LAYER M3 ;
        RECT 20.93 7.56 21.21 13.86 ;
  LAYER M1 ;
        RECT 23.525 7.055 23.775 7.225 ;
  LAYER M2 ;
        RECT 23.48 7 23.82 7.28 ;
  LAYER M1 ;
        RECT 23.525 7.475 23.775 7.645 ;
  LAYER M2 ;
        RECT 23.48 7.42 23.82 7.7 ;
  LAYER M2 ;
        RECT 11.88 7.42 12.2 7.7 ;
  LAYER M3 ;
        RECT 11.9 7.4 12.18 7.72 ;
  LAYER M1 ;
        RECT 23.525 7.055 23.775 7.225 ;
  LAYER M2 ;
        RECT 23.48 7 23.82 7.28 ;
  LAYER M1 ;
        RECT 23.525 7.475 23.775 7.645 ;
  LAYER M2 ;
        RECT 23.48 7.42 23.82 7.7 ;
  LAYER M2 ;
        RECT 11.88 7.42 12.2 7.7 ;
  LAYER M3 ;
        RECT 11.9 7.4 12.18 7.72 ;
  LAYER M1 ;
        RECT 23.525 7.055 23.775 7.225 ;
  LAYER M2 ;
        RECT 23.48 7 23.82 7.28 ;
  LAYER M1 ;
        RECT 23.525 7.475 23.775 7.645 ;
  LAYER M2 ;
        RECT 23.48 7.42 23.82 7.7 ;
  LAYER M2 ;
        RECT 11.88 7.42 12.2 7.7 ;
  LAYER M3 ;
        RECT 11.9 7.4 12.18 7.72 ;
  LAYER M2 ;
        RECT 20.91 7.42 21.23 7.7 ;
  LAYER M3 ;
        RECT 20.93 7.4 21.21 7.72 ;
  LAYER M1 ;
        RECT 23.525 7.055 23.775 7.225 ;
  LAYER M2 ;
        RECT 23.48 7 23.82 7.28 ;
  LAYER M1 ;
        RECT 23.525 7.475 23.775 7.645 ;
  LAYER M2 ;
        RECT 23.48 7.42 23.82 7.7 ;
  LAYER M2 ;
        RECT 11.88 7.42 12.2 7.7 ;
  LAYER M3 ;
        RECT 11.9 7.4 12.18 7.72 ;
  LAYER M2 ;
        RECT 20.91 7.42 21.23 7.7 ;
  LAYER M3 ;
        RECT 20.93 7.4 21.21 7.72 ;
  LAYER M2 ;
        RECT 27.78 7 28.98 7.28 ;
  LAYER M3 ;
        RECT 32.11 13.7 32.39 18.22 ;
  LAYER M3 ;
        RECT 41.14 2.78 41.42 8.98 ;
  LAYER M2 ;
        RECT 28.81 7 29.67 7.28 ;
  LAYER M3 ;
        RECT 29.53 7.14 29.81 9.66 ;
  LAYER M2 ;
        RECT 29.67 9.52 32.25 9.8 ;
  LAYER M3 ;
        RECT 32.11 9.66 32.39 13.86 ;
  LAYER M2 ;
        RECT 32.25 9.52 41.28 9.8 ;
  LAYER M3 ;
        RECT 41.14 8.82 41.42 9.66 ;
  LAYER M2 ;
        RECT 29.51 7 29.83 7.28 ;
  LAYER M3 ;
        RECT 29.53 6.98 29.81 7.3 ;
  LAYER M2 ;
        RECT 29.51 9.52 29.83 9.8 ;
  LAYER M3 ;
        RECT 29.53 9.5 29.81 9.82 ;
  LAYER M2 ;
        RECT 32.09 9.52 32.41 9.8 ;
  LAYER M3 ;
        RECT 32.11 9.5 32.39 9.82 ;
  LAYER M2 ;
        RECT 29.51 7 29.83 7.28 ;
  LAYER M3 ;
        RECT 29.53 6.98 29.81 7.3 ;
  LAYER M2 ;
        RECT 29.51 9.52 29.83 9.8 ;
  LAYER M3 ;
        RECT 29.53 9.5 29.81 9.82 ;
  LAYER M2 ;
        RECT 32.09 9.52 32.41 9.8 ;
  LAYER M3 ;
        RECT 32.11 9.5 32.39 9.82 ;
  LAYER M2 ;
        RECT 29.51 7 29.83 7.28 ;
  LAYER M3 ;
        RECT 29.53 6.98 29.81 7.3 ;
  LAYER M2 ;
        RECT 29.51 9.52 29.83 9.8 ;
  LAYER M3 ;
        RECT 29.53 9.5 29.81 9.82 ;
  LAYER M2 ;
        RECT 32.09 9.52 32.41 9.8 ;
  LAYER M3 ;
        RECT 32.11 9.5 32.39 9.82 ;
  LAYER M2 ;
        RECT 41.12 9.52 41.44 9.8 ;
  LAYER M3 ;
        RECT 41.14 9.5 41.42 9.82 ;
  LAYER M2 ;
        RECT 29.51 7 29.83 7.28 ;
  LAYER M3 ;
        RECT 29.53 6.98 29.81 7.3 ;
  LAYER M2 ;
        RECT 29.51 9.52 29.83 9.8 ;
  LAYER M3 ;
        RECT 29.53 9.5 29.81 9.82 ;
  LAYER M2 ;
        RECT 32.09 9.52 32.41 9.8 ;
  LAYER M3 ;
        RECT 32.11 9.5 32.39 9.82 ;
  LAYER M2 ;
        RECT 41.12 9.52 41.44 9.8 ;
  LAYER M3 ;
        RECT 41.14 9.5 41.42 9.82 ;
  LAYER M2 ;
        RECT 24.77 6.58 25.97 6.86 ;
  LAYER M2 ;
        RECT 27.35 6.58 28.55 6.86 ;
  LAYER M2 ;
        RECT 26.92 7.84 28.12 8.12 ;
  LAYER M2 ;
        RECT 25.8 6.58 27.52 6.86 ;
  LAYER M2 ;
        RECT 26.93 6.58 27.25 6.86 ;
  LAYER M1 ;
        RECT 26.965 6.72 27.215 7.98 ;
  LAYER M2 ;
        RECT 26.93 7.84 27.25 8.12 ;
  LAYER M1 ;
        RECT 26.965 6.635 27.215 6.805 ;
  LAYER M2 ;
        RECT 26.92 6.58 27.26 6.86 ;
  LAYER M1 ;
        RECT 26.965 7.895 27.215 8.065 ;
  LAYER M2 ;
        RECT 26.92 7.84 27.26 8.12 ;
  LAYER M1 ;
        RECT 26.965 6.635 27.215 6.805 ;
  LAYER M2 ;
        RECT 26.92 6.58 27.26 6.86 ;
  LAYER M1 ;
        RECT 26.965 7.895 27.215 8.065 ;
  LAYER M2 ;
        RECT 26.92 7.84 27.26 8.12 ;
  LAYER M1 ;
        RECT 25.245 7.895 25.495 11.425 ;
  LAYER M1 ;
        RECT 25.245 11.675 25.495 12.685 ;
  LAYER M1 ;
        RECT 25.245 13.775 25.495 14.785 ;
  LAYER M1 ;
        RECT 25.675 7.895 25.925 11.425 ;
  LAYER M1 ;
        RECT 24.815 7.895 25.065 11.425 ;
  LAYER M2 ;
        RECT 25.2 7.84 26.4 8.12 ;
  LAYER M2 ;
        RECT 25.2 12.04 26.4 12.32 ;
  LAYER M2 ;
        RECT 24.77 8.26 25.97 8.54 ;
  LAYER M2 ;
        RECT 24.77 14.14 25.97 14.42 ;
  LAYER M3 ;
        RECT 25.23 7.82 25.51 12.34 ;
  LAYER M3 ;
        RECT 24.8 8.24 25.08 14.44 ;
  LAYER M1 ;
        RECT 36.425 13.775 36.675 17.305 ;
  LAYER M1 ;
        RECT 36.425 17.555 36.675 18.565 ;
  LAYER M1 ;
        RECT 36.425 19.655 36.675 20.665 ;
  LAYER M1 ;
        RECT 35.995 13.775 36.245 17.305 ;
  LAYER M1 ;
        RECT 36.855 13.775 37.105 17.305 ;
  LAYER M1 ;
        RECT 37.285 13.775 37.535 17.305 ;
  LAYER M1 ;
        RECT 37.285 17.555 37.535 18.565 ;
  LAYER M1 ;
        RECT 37.285 19.655 37.535 20.665 ;
  LAYER M1 ;
        RECT 37.715 13.775 37.965 17.305 ;
  LAYER M1 ;
        RECT 38.145 13.775 38.395 17.305 ;
  LAYER M1 ;
        RECT 38.145 17.555 38.395 18.565 ;
  LAYER M1 ;
        RECT 38.145 19.655 38.395 20.665 ;
  LAYER M1 ;
        RECT 38.575 13.775 38.825 17.305 ;
  LAYER M1 ;
        RECT 39.005 13.775 39.255 17.305 ;
  LAYER M1 ;
        RECT 39.005 17.555 39.255 18.565 ;
  LAYER M1 ;
        RECT 39.005 19.655 39.255 20.665 ;
  LAYER M1 ;
        RECT 39.435 13.775 39.685 17.305 ;
  LAYER M1 ;
        RECT 39.865 13.775 40.115 17.305 ;
  LAYER M1 ;
        RECT 39.865 17.555 40.115 18.565 ;
  LAYER M1 ;
        RECT 39.865 19.655 40.115 20.665 ;
  LAYER M1 ;
        RECT 40.295 13.775 40.545 17.305 ;
  LAYER M1 ;
        RECT 40.725 13.775 40.975 17.305 ;
  LAYER M1 ;
        RECT 40.725 17.555 40.975 18.565 ;
  LAYER M1 ;
        RECT 40.725 19.655 40.975 20.665 ;
  LAYER M1 ;
        RECT 41.155 13.775 41.405 17.305 ;
  LAYER M1 ;
        RECT 41.585 13.775 41.835 17.305 ;
  LAYER M1 ;
        RECT 41.585 17.555 41.835 18.565 ;
  LAYER M1 ;
        RECT 41.585 19.655 41.835 20.665 ;
  LAYER M1 ;
        RECT 42.015 13.775 42.265 17.305 ;
  LAYER M1 ;
        RECT 42.445 13.775 42.695 17.305 ;
  LAYER M1 ;
        RECT 42.445 17.555 42.695 18.565 ;
  LAYER M1 ;
        RECT 42.445 19.655 42.695 20.665 ;
  LAYER M1 ;
        RECT 42.875 13.775 43.125 17.305 ;
  LAYER M1 ;
        RECT 43.305 13.775 43.555 17.305 ;
  LAYER M1 ;
        RECT 43.305 17.555 43.555 18.565 ;
  LAYER M1 ;
        RECT 43.305 19.655 43.555 20.665 ;
  LAYER M1 ;
        RECT 43.735 13.775 43.985 17.305 ;
  LAYER M1 ;
        RECT 44.165 13.775 44.415 17.305 ;
  LAYER M1 ;
        RECT 44.165 17.555 44.415 18.565 ;
  LAYER M1 ;
        RECT 44.165 19.655 44.415 20.665 ;
  LAYER M1 ;
        RECT 44.595 13.775 44.845 17.305 ;
  LAYER M1 ;
        RECT 45.025 13.775 45.275 17.305 ;
  LAYER M1 ;
        RECT 45.025 17.555 45.275 18.565 ;
  LAYER M1 ;
        RECT 45.025 19.655 45.275 20.665 ;
  LAYER M1 ;
        RECT 45.455 13.775 45.705 17.305 ;
  LAYER M1 ;
        RECT 45.885 13.775 46.135 17.305 ;
  LAYER M1 ;
        RECT 45.885 17.555 46.135 18.565 ;
  LAYER M1 ;
        RECT 45.885 19.655 46.135 20.665 ;
  LAYER M1 ;
        RECT 46.315 13.775 46.565 17.305 ;
  LAYER M1 ;
        RECT 46.745 13.775 46.995 17.305 ;
  LAYER M1 ;
        RECT 46.745 17.555 46.995 18.565 ;
  LAYER M1 ;
        RECT 46.745 19.655 46.995 20.665 ;
  LAYER M1 ;
        RECT 47.175 13.775 47.425 17.305 ;
  LAYER M1 ;
        RECT 47.605 13.775 47.855 17.305 ;
  LAYER M1 ;
        RECT 47.605 17.555 47.855 18.565 ;
  LAYER M1 ;
        RECT 47.605 19.655 47.855 20.665 ;
  LAYER M1 ;
        RECT 48.035 13.775 48.285 17.305 ;
  LAYER M2 ;
        RECT 36.38 13.72 47.9 14 ;
  LAYER M2 ;
        RECT 36.38 17.92 47.9 18.2 ;
  LAYER M2 ;
        RECT 35.95 14.14 48.33 14.42 ;
  LAYER M2 ;
        RECT 36.38 20.02 47.9 20.3 ;
  LAYER M3 ;
        RECT 42 13.7 42.28 18.22 ;
  LAYER M3 ;
        RECT 42.43 14.12 42.71 20.32 ;
  LAYER M1 ;
        RECT 22.665 13.775 22.915 17.305 ;
  LAYER M1 ;
        RECT 22.665 17.555 22.915 18.565 ;
  LAYER M1 ;
        RECT 22.665 19.655 22.915 20.665 ;
  LAYER M1 ;
        RECT 23.095 13.775 23.345 17.305 ;
  LAYER M1 ;
        RECT 22.235 13.775 22.485 17.305 ;
  LAYER M1 ;
        RECT 21.805 13.775 22.055 17.305 ;
  LAYER M1 ;
        RECT 21.805 17.555 22.055 18.565 ;
  LAYER M1 ;
        RECT 21.805 19.655 22.055 20.665 ;
  LAYER M1 ;
        RECT 21.375 13.775 21.625 17.305 ;
  LAYER M1 ;
        RECT 20.945 13.775 21.195 17.305 ;
  LAYER M1 ;
        RECT 20.945 17.555 21.195 18.565 ;
  LAYER M1 ;
        RECT 20.945 19.655 21.195 20.665 ;
  LAYER M1 ;
        RECT 20.515 13.775 20.765 17.305 ;
  LAYER M1 ;
        RECT 20.085 13.775 20.335 17.305 ;
  LAYER M1 ;
        RECT 20.085 17.555 20.335 18.565 ;
  LAYER M1 ;
        RECT 20.085 19.655 20.335 20.665 ;
  LAYER M1 ;
        RECT 19.655 13.775 19.905 17.305 ;
  LAYER M1 ;
        RECT 19.225 13.775 19.475 17.305 ;
  LAYER M1 ;
        RECT 19.225 17.555 19.475 18.565 ;
  LAYER M1 ;
        RECT 19.225 19.655 19.475 20.665 ;
  LAYER M1 ;
        RECT 18.795 13.775 19.045 17.305 ;
  LAYER M2 ;
        RECT 19.18 13.72 22.96 14 ;
  LAYER M2 ;
        RECT 19.18 17.92 22.96 18.2 ;
  LAYER M2 ;
        RECT 19.18 20.02 22.96 20.3 ;
  LAYER M2 ;
        RECT 18.75 14.14 23.39 14.42 ;
  LAYER M3 ;
        RECT 20.93 13.7 21.21 18.22 ;
  LAYER M3 ;
        RECT 20.5 14.12 20.78 20.32 ;
  LAYER M1 ;
        RECT 30.405 13.775 30.655 17.305 ;
  LAYER M1 ;
        RECT 30.405 17.555 30.655 18.565 ;
  LAYER M1 ;
        RECT 30.405 19.655 30.655 20.665 ;
  LAYER M1 ;
        RECT 29.975 13.775 30.225 17.305 ;
  LAYER M1 ;
        RECT 30.835 13.775 31.085 17.305 ;
  LAYER M1 ;
        RECT 31.265 13.775 31.515 17.305 ;
  LAYER M1 ;
        RECT 31.265 17.555 31.515 18.565 ;
  LAYER M1 ;
        RECT 31.265 19.655 31.515 20.665 ;
  LAYER M1 ;
        RECT 31.695 13.775 31.945 17.305 ;
  LAYER M1 ;
        RECT 32.125 13.775 32.375 17.305 ;
  LAYER M1 ;
        RECT 32.125 17.555 32.375 18.565 ;
  LAYER M1 ;
        RECT 32.125 19.655 32.375 20.665 ;
  LAYER M1 ;
        RECT 32.555 13.775 32.805 17.305 ;
  LAYER M1 ;
        RECT 32.985 13.775 33.235 17.305 ;
  LAYER M1 ;
        RECT 32.985 17.555 33.235 18.565 ;
  LAYER M1 ;
        RECT 32.985 19.655 33.235 20.665 ;
  LAYER M1 ;
        RECT 33.415 13.775 33.665 17.305 ;
  LAYER M1 ;
        RECT 33.845 13.775 34.095 17.305 ;
  LAYER M1 ;
        RECT 33.845 17.555 34.095 18.565 ;
  LAYER M1 ;
        RECT 33.845 19.655 34.095 20.665 ;
  LAYER M1 ;
        RECT 34.275 13.775 34.525 17.305 ;
  LAYER M2 ;
        RECT 30.36 13.72 34.14 14 ;
  LAYER M2 ;
        RECT 30.36 17.92 34.14 18.2 ;
  LAYER M2 ;
        RECT 30.36 20.02 34.14 20.3 ;
  LAYER M2 ;
        RECT 29.93 14.14 34.57 14.42 ;
  LAYER M3 ;
        RECT 32.11 13.7 32.39 18.22 ;
  LAYER M3 ;
        RECT 32.54 14.12 32.82 20.32 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 17.305 ;
  LAYER M1 ;
        RECT 16.645 17.555 16.895 18.565 ;
  LAYER M1 ;
        RECT 16.645 19.655 16.895 20.665 ;
  LAYER M1 ;
        RECT 17.075 13.775 17.325 17.305 ;
  LAYER M1 ;
        RECT 16.215 13.775 16.465 17.305 ;
  LAYER M1 ;
        RECT 15.785 13.775 16.035 17.305 ;
  LAYER M1 ;
        RECT 15.785 17.555 16.035 18.565 ;
  LAYER M1 ;
        RECT 15.785 19.655 16.035 20.665 ;
  LAYER M1 ;
        RECT 15.355 13.775 15.605 17.305 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 17.305 ;
  LAYER M1 ;
        RECT 14.925 17.555 15.175 18.565 ;
  LAYER M1 ;
        RECT 14.925 19.655 15.175 20.665 ;
  LAYER M1 ;
        RECT 14.495 13.775 14.745 17.305 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 17.305 ;
  LAYER M1 ;
        RECT 14.065 17.555 14.315 18.565 ;
  LAYER M1 ;
        RECT 14.065 19.655 14.315 20.665 ;
  LAYER M1 ;
        RECT 13.635 13.775 13.885 17.305 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 17.305 ;
  LAYER M1 ;
        RECT 13.205 17.555 13.455 18.565 ;
  LAYER M1 ;
        RECT 13.205 19.655 13.455 20.665 ;
  LAYER M1 ;
        RECT 12.775 13.775 13.025 17.305 ;
  LAYER M1 ;
        RECT 12.345 13.775 12.595 17.305 ;
  LAYER M1 ;
        RECT 12.345 17.555 12.595 18.565 ;
  LAYER M1 ;
        RECT 12.345 19.655 12.595 20.665 ;
  LAYER M1 ;
        RECT 11.915 13.775 12.165 17.305 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 17.305 ;
  LAYER M1 ;
        RECT 11.485 17.555 11.735 18.565 ;
  LAYER M1 ;
        RECT 11.485 19.655 11.735 20.665 ;
  LAYER M1 ;
        RECT 11.055 13.775 11.305 17.305 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 17.305 ;
  LAYER M1 ;
        RECT 10.625 17.555 10.875 18.565 ;
  LAYER M1 ;
        RECT 10.625 19.655 10.875 20.665 ;
  LAYER M1 ;
        RECT 10.195 13.775 10.445 17.305 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 17.305 ;
  LAYER M1 ;
        RECT 9.765 17.555 10.015 18.565 ;
  LAYER M1 ;
        RECT 9.765 19.655 10.015 20.665 ;
  LAYER M1 ;
        RECT 9.335 13.775 9.585 17.305 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 17.305 ;
  LAYER M1 ;
        RECT 8.905 17.555 9.155 18.565 ;
  LAYER M1 ;
        RECT 8.905 19.655 9.155 20.665 ;
  LAYER M1 ;
        RECT 8.475 13.775 8.725 17.305 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 17.305 ;
  LAYER M1 ;
        RECT 8.045 17.555 8.295 18.565 ;
  LAYER M1 ;
        RECT 8.045 19.655 8.295 20.665 ;
  LAYER M1 ;
        RECT 7.615 13.775 7.865 17.305 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 17.305 ;
  LAYER M1 ;
        RECT 7.185 17.555 7.435 18.565 ;
  LAYER M1 ;
        RECT 7.185 19.655 7.435 20.665 ;
  LAYER M1 ;
        RECT 6.755 13.775 7.005 17.305 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 17.305 ;
  LAYER M1 ;
        RECT 6.325 17.555 6.575 18.565 ;
  LAYER M1 ;
        RECT 6.325 19.655 6.575 20.665 ;
  LAYER M1 ;
        RECT 5.895 13.775 6.145 17.305 ;
  LAYER M1 ;
        RECT 5.465 13.775 5.715 17.305 ;
  LAYER M1 ;
        RECT 5.465 17.555 5.715 18.565 ;
  LAYER M1 ;
        RECT 5.465 19.655 5.715 20.665 ;
  LAYER M1 ;
        RECT 5.035 13.775 5.285 17.305 ;
  LAYER M2 ;
        RECT 4.99 14.14 17.37 14.42 ;
  LAYER M2 ;
        RECT 5.42 20.02 16.94 20.3 ;
  LAYER M2 ;
        RECT 5.42 13.72 16.94 14 ;
  LAYER M2 ;
        RECT 5.42 17.92 16.94 18.2 ;
  LAYER M3 ;
        RECT 10.61 14.12 10.89 20.32 ;
  LAYER M1 ;
        RECT 27.825 7.895 28.075 11.425 ;
  LAYER M1 ;
        RECT 27.825 11.675 28.075 12.685 ;
  LAYER M1 ;
        RECT 27.825 13.775 28.075 14.785 ;
  LAYER M1 ;
        RECT 27.395 7.895 27.645 11.425 ;
  LAYER M1 ;
        RECT 28.255 7.895 28.505 11.425 ;
  LAYER M2 ;
        RECT 27.35 8.26 28.55 8.54 ;
  LAYER M2 ;
        RECT 27.35 14.14 28.55 14.42 ;
  LAYER M2 ;
        RECT 26.92 7.84 28.12 8.12 ;
  LAYER M2 ;
        RECT 26.92 12.04 28.12 12.32 ;
  LAYER M3 ;
        RECT 28.24 8.24 28.52 14.44 ;
  LAYER M1 ;
        RECT 30.405 9.575 30.655 13.105 ;
  LAYER M1 ;
        RECT 30.405 8.315 30.655 9.325 ;
  LAYER M1 ;
        RECT 30.405 3.695 30.655 7.225 ;
  LAYER M1 ;
        RECT 30.405 2.435 30.655 3.445 ;
  LAYER M1 ;
        RECT 30.405 0.335 30.655 1.345 ;
  LAYER M1 ;
        RECT 29.975 9.575 30.225 13.105 ;
  LAYER M1 ;
        RECT 29.975 3.695 30.225 7.225 ;
  LAYER M1 ;
        RECT 30.835 9.575 31.085 13.105 ;
  LAYER M1 ;
        RECT 30.835 3.695 31.085 7.225 ;
  LAYER M1 ;
        RECT 31.265 9.575 31.515 13.105 ;
  LAYER M1 ;
        RECT 31.265 8.315 31.515 9.325 ;
  LAYER M1 ;
        RECT 31.265 3.695 31.515 7.225 ;
  LAYER M1 ;
        RECT 31.265 2.435 31.515 3.445 ;
  LAYER M1 ;
        RECT 31.265 0.335 31.515 1.345 ;
  LAYER M1 ;
        RECT 31.695 9.575 31.945 13.105 ;
  LAYER M1 ;
        RECT 31.695 3.695 31.945 7.225 ;
  LAYER M1 ;
        RECT 32.125 9.575 32.375 13.105 ;
  LAYER M1 ;
        RECT 32.125 8.315 32.375 9.325 ;
  LAYER M1 ;
        RECT 32.125 3.695 32.375 7.225 ;
  LAYER M1 ;
        RECT 32.125 2.435 32.375 3.445 ;
  LAYER M1 ;
        RECT 32.125 0.335 32.375 1.345 ;
  LAYER M1 ;
        RECT 32.555 9.575 32.805 13.105 ;
  LAYER M1 ;
        RECT 32.555 3.695 32.805 7.225 ;
  LAYER M1 ;
        RECT 32.985 9.575 33.235 13.105 ;
  LAYER M1 ;
        RECT 32.985 8.315 33.235 9.325 ;
  LAYER M1 ;
        RECT 32.985 3.695 33.235 7.225 ;
  LAYER M1 ;
        RECT 32.985 2.435 33.235 3.445 ;
  LAYER M1 ;
        RECT 32.985 0.335 33.235 1.345 ;
  LAYER M1 ;
        RECT 33.415 9.575 33.665 13.105 ;
  LAYER M1 ;
        RECT 33.415 3.695 33.665 7.225 ;
  LAYER M1 ;
        RECT 33.845 9.575 34.095 13.105 ;
  LAYER M1 ;
        RECT 33.845 8.315 34.095 9.325 ;
  LAYER M1 ;
        RECT 33.845 3.695 34.095 7.225 ;
  LAYER M1 ;
        RECT 33.845 2.435 34.095 3.445 ;
  LAYER M1 ;
        RECT 33.845 0.335 34.095 1.345 ;
  LAYER M1 ;
        RECT 34.275 9.575 34.525 13.105 ;
  LAYER M1 ;
        RECT 34.275 3.695 34.525 7.225 ;
  LAYER M1 ;
        RECT 34.705 9.575 34.955 13.105 ;
  LAYER M1 ;
        RECT 34.705 8.315 34.955 9.325 ;
  LAYER M1 ;
        RECT 34.705 3.695 34.955 7.225 ;
  LAYER M1 ;
        RECT 34.705 2.435 34.955 3.445 ;
  LAYER M1 ;
        RECT 34.705 0.335 34.955 1.345 ;
  LAYER M1 ;
        RECT 35.135 9.575 35.385 13.105 ;
  LAYER M1 ;
        RECT 35.135 3.695 35.385 7.225 ;
  LAYER M1 ;
        RECT 35.565 9.575 35.815 13.105 ;
  LAYER M1 ;
        RECT 35.565 8.315 35.815 9.325 ;
  LAYER M1 ;
        RECT 35.565 3.695 35.815 7.225 ;
  LAYER M1 ;
        RECT 35.565 2.435 35.815 3.445 ;
  LAYER M1 ;
        RECT 35.565 0.335 35.815 1.345 ;
  LAYER M1 ;
        RECT 35.995 9.575 36.245 13.105 ;
  LAYER M1 ;
        RECT 35.995 3.695 36.245 7.225 ;
  LAYER M1 ;
        RECT 36.425 9.575 36.675 13.105 ;
  LAYER M1 ;
        RECT 36.425 8.315 36.675 9.325 ;
  LAYER M1 ;
        RECT 36.425 3.695 36.675 7.225 ;
  LAYER M1 ;
        RECT 36.425 2.435 36.675 3.445 ;
  LAYER M1 ;
        RECT 36.425 0.335 36.675 1.345 ;
  LAYER M1 ;
        RECT 36.855 9.575 37.105 13.105 ;
  LAYER M1 ;
        RECT 36.855 3.695 37.105 7.225 ;
  LAYER M1 ;
        RECT 37.285 9.575 37.535 13.105 ;
  LAYER M1 ;
        RECT 37.285 8.315 37.535 9.325 ;
  LAYER M1 ;
        RECT 37.285 3.695 37.535 7.225 ;
  LAYER M1 ;
        RECT 37.285 2.435 37.535 3.445 ;
  LAYER M1 ;
        RECT 37.285 0.335 37.535 1.345 ;
  LAYER M1 ;
        RECT 37.715 9.575 37.965 13.105 ;
  LAYER M1 ;
        RECT 37.715 3.695 37.965 7.225 ;
  LAYER M1 ;
        RECT 38.145 9.575 38.395 13.105 ;
  LAYER M1 ;
        RECT 38.145 8.315 38.395 9.325 ;
  LAYER M1 ;
        RECT 38.145 3.695 38.395 7.225 ;
  LAYER M1 ;
        RECT 38.145 2.435 38.395 3.445 ;
  LAYER M1 ;
        RECT 38.145 0.335 38.395 1.345 ;
  LAYER M1 ;
        RECT 38.575 9.575 38.825 13.105 ;
  LAYER M1 ;
        RECT 38.575 3.695 38.825 7.225 ;
  LAYER M1 ;
        RECT 39.005 9.575 39.255 13.105 ;
  LAYER M1 ;
        RECT 39.005 8.315 39.255 9.325 ;
  LAYER M1 ;
        RECT 39.005 3.695 39.255 7.225 ;
  LAYER M1 ;
        RECT 39.005 2.435 39.255 3.445 ;
  LAYER M1 ;
        RECT 39.005 0.335 39.255 1.345 ;
  LAYER M1 ;
        RECT 39.435 9.575 39.685 13.105 ;
  LAYER M1 ;
        RECT 39.435 3.695 39.685 7.225 ;
  LAYER M1 ;
        RECT 39.865 9.575 40.115 13.105 ;
  LAYER M1 ;
        RECT 39.865 8.315 40.115 9.325 ;
  LAYER M1 ;
        RECT 39.865 3.695 40.115 7.225 ;
  LAYER M1 ;
        RECT 39.865 2.435 40.115 3.445 ;
  LAYER M1 ;
        RECT 39.865 0.335 40.115 1.345 ;
  LAYER M1 ;
        RECT 40.295 9.575 40.545 13.105 ;
  LAYER M1 ;
        RECT 40.295 3.695 40.545 7.225 ;
  LAYER M1 ;
        RECT 40.725 9.575 40.975 13.105 ;
  LAYER M1 ;
        RECT 40.725 8.315 40.975 9.325 ;
  LAYER M1 ;
        RECT 40.725 3.695 40.975 7.225 ;
  LAYER M1 ;
        RECT 40.725 2.435 40.975 3.445 ;
  LAYER M1 ;
        RECT 40.725 0.335 40.975 1.345 ;
  LAYER M1 ;
        RECT 41.155 9.575 41.405 13.105 ;
  LAYER M1 ;
        RECT 41.155 3.695 41.405 7.225 ;
  LAYER M1 ;
        RECT 41.585 9.575 41.835 13.105 ;
  LAYER M1 ;
        RECT 41.585 8.315 41.835 9.325 ;
  LAYER M1 ;
        RECT 41.585 3.695 41.835 7.225 ;
  LAYER M1 ;
        RECT 41.585 2.435 41.835 3.445 ;
  LAYER M1 ;
        RECT 41.585 0.335 41.835 1.345 ;
  LAYER M1 ;
        RECT 42.015 9.575 42.265 13.105 ;
  LAYER M1 ;
        RECT 42.015 3.695 42.265 7.225 ;
  LAYER M1 ;
        RECT 42.445 9.575 42.695 13.105 ;
  LAYER M1 ;
        RECT 42.445 8.315 42.695 9.325 ;
  LAYER M1 ;
        RECT 42.445 3.695 42.695 7.225 ;
  LAYER M1 ;
        RECT 42.445 2.435 42.695 3.445 ;
  LAYER M1 ;
        RECT 42.445 0.335 42.695 1.345 ;
  LAYER M1 ;
        RECT 42.875 9.575 43.125 13.105 ;
  LAYER M1 ;
        RECT 42.875 3.695 43.125 7.225 ;
  LAYER M1 ;
        RECT 43.305 9.575 43.555 13.105 ;
  LAYER M1 ;
        RECT 43.305 8.315 43.555 9.325 ;
  LAYER M1 ;
        RECT 43.305 3.695 43.555 7.225 ;
  LAYER M1 ;
        RECT 43.305 2.435 43.555 3.445 ;
  LAYER M1 ;
        RECT 43.305 0.335 43.555 1.345 ;
  LAYER M1 ;
        RECT 43.735 9.575 43.985 13.105 ;
  LAYER M1 ;
        RECT 43.735 3.695 43.985 7.225 ;
  LAYER M1 ;
        RECT 44.165 9.575 44.415 13.105 ;
  LAYER M1 ;
        RECT 44.165 8.315 44.415 9.325 ;
  LAYER M1 ;
        RECT 44.165 3.695 44.415 7.225 ;
  LAYER M1 ;
        RECT 44.165 2.435 44.415 3.445 ;
  LAYER M1 ;
        RECT 44.165 0.335 44.415 1.345 ;
  LAYER M1 ;
        RECT 44.595 9.575 44.845 13.105 ;
  LAYER M1 ;
        RECT 44.595 3.695 44.845 7.225 ;
  LAYER M1 ;
        RECT 45.025 9.575 45.275 13.105 ;
  LAYER M1 ;
        RECT 45.025 8.315 45.275 9.325 ;
  LAYER M1 ;
        RECT 45.025 3.695 45.275 7.225 ;
  LAYER M1 ;
        RECT 45.025 2.435 45.275 3.445 ;
  LAYER M1 ;
        RECT 45.025 0.335 45.275 1.345 ;
  LAYER M1 ;
        RECT 45.455 9.575 45.705 13.105 ;
  LAYER M1 ;
        RECT 45.455 3.695 45.705 7.225 ;
  LAYER M1 ;
        RECT 45.885 9.575 46.135 13.105 ;
  LAYER M1 ;
        RECT 45.885 8.315 46.135 9.325 ;
  LAYER M1 ;
        RECT 45.885 3.695 46.135 7.225 ;
  LAYER M1 ;
        RECT 45.885 2.435 46.135 3.445 ;
  LAYER M1 ;
        RECT 45.885 0.335 46.135 1.345 ;
  LAYER M1 ;
        RECT 46.315 9.575 46.565 13.105 ;
  LAYER M1 ;
        RECT 46.315 3.695 46.565 7.225 ;
  LAYER M1 ;
        RECT 46.745 9.575 46.995 13.105 ;
  LAYER M1 ;
        RECT 46.745 8.315 46.995 9.325 ;
  LAYER M1 ;
        RECT 46.745 3.695 46.995 7.225 ;
  LAYER M1 ;
        RECT 46.745 2.435 46.995 3.445 ;
  LAYER M1 ;
        RECT 46.745 0.335 46.995 1.345 ;
  LAYER M1 ;
        RECT 47.175 9.575 47.425 13.105 ;
  LAYER M1 ;
        RECT 47.175 3.695 47.425 7.225 ;
  LAYER M1 ;
        RECT 47.605 9.575 47.855 13.105 ;
  LAYER M1 ;
        RECT 47.605 8.315 47.855 9.325 ;
  LAYER M1 ;
        RECT 47.605 3.695 47.855 7.225 ;
  LAYER M1 ;
        RECT 47.605 2.435 47.855 3.445 ;
  LAYER M1 ;
        RECT 47.605 0.335 47.855 1.345 ;
  LAYER M1 ;
        RECT 48.035 9.575 48.285 13.105 ;
  LAYER M1 ;
        RECT 48.035 3.695 48.285 7.225 ;
  LAYER M1 ;
        RECT 48.465 9.575 48.715 13.105 ;
  LAYER M1 ;
        RECT 48.465 8.315 48.715 9.325 ;
  LAYER M1 ;
        RECT 48.465 3.695 48.715 7.225 ;
  LAYER M1 ;
        RECT 48.465 2.435 48.715 3.445 ;
  LAYER M1 ;
        RECT 48.465 0.335 48.715 1.345 ;
  LAYER M1 ;
        RECT 48.895 9.575 49.145 13.105 ;
  LAYER M1 ;
        RECT 48.895 3.695 49.145 7.225 ;
  LAYER M1 ;
        RECT 49.325 9.575 49.575 13.105 ;
  LAYER M1 ;
        RECT 49.325 8.315 49.575 9.325 ;
  LAYER M1 ;
        RECT 49.325 3.695 49.575 7.225 ;
  LAYER M1 ;
        RECT 49.325 2.435 49.575 3.445 ;
  LAYER M1 ;
        RECT 49.325 0.335 49.575 1.345 ;
  LAYER M1 ;
        RECT 49.755 9.575 50.005 13.105 ;
  LAYER M1 ;
        RECT 49.755 3.695 50.005 7.225 ;
  LAYER M1 ;
        RECT 50.185 9.575 50.435 13.105 ;
  LAYER M1 ;
        RECT 50.185 8.315 50.435 9.325 ;
  LAYER M1 ;
        RECT 50.185 3.695 50.435 7.225 ;
  LAYER M1 ;
        RECT 50.185 2.435 50.435 3.445 ;
  LAYER M1 ;
        RECT 50.185 0.335 50.435 1.345 ;
  LAYER M1 ;
        RECT 50.615 9.575 50.865 13.105 ;
  LAYER M1 ;
        RECT 50.615 3.695 50.865 7.225 ;
  LAYER M1 ;
        RECT 51.045 9.575 51.295 13.105 ;
  LAYER M1 ;
        RECT 51.045 8.315 51.295 9.325 ;
  LAYER M1 ;
        RECT 51.045 3.695 51.295 7.225 ;
  LAYER M1 ;
        RECT 51.045 2.435 51.295 3.445 ;
  LAYER M1 ;
        RECT 51.045 0.335 51.295 1.345 ;
  LAYER M1 ;
        RECT 51.475 9.575 51.725 13.105 ;
  LAYER M1 ;
        RECT 51.475 3.695 51.725 7.225 ;
  LAYER M1 ;
        RECT 51.905 9.575 52.155 13.105 ;
  LAYER M1 ;
        RECT 51.905 8.315 52.155 9.325 ;
  LAYER M1 ;
        RECT 51.905 3.695 52.155 7.225 ;
  LAYER M1 ;
        RECT 51.905 2.435 52.155 3.445 ;
  LAYER M1 ;
        RECT 51.905 0.335 52.155 1.345 ;
  LAYER M1 ;
        RECT 52.335 9.575 52.585 13.105 ;
  LAYER M1 ;
        RECT 52.335 3.695 52.585 7.225 ;
  LAYER M2 ;
        RECT 30.36 12.88 52.2 13.16 ;
  LAYER M2 ;
        RECT 30.36 8.68 52.2 8.96 ;
  LAYER M2 ;
        RECT 29.93 12.46 52.63 12.74 ;
  LAYER M2 ;
        RECT 30.36 7 52.2 7.28 ;
  LAYER M2 ;
        RECT 30.36 2.8 52.2 3.08 ;
  LAYER M2 ;
        RECT 29.93 6.58 52.63 6.86 ;
  LAYER M2 ;
        RECT 30.36 0.7 52.2 0.98 ;
  LAYER M3 ;
        RECT 40.71 6.98 40.99 13.18 ;
  LAYER M3 ;
        RECT 41.14 2.78 41.42 8.98 ;
  LAYER M3 ;
        RECT 41.57 0.68 41.85 12.76 ;
  LAYER M1 ;
        RECT 22.665 9.575 22.915 13.105 ;
  LAYER M1 ;
        RECT 22.665 8.315 22.915 9.325 ;
  LAYER M1 ;
        RECT 22.665 3.695 22.915 7.225 ;
  LAYER M1 ;
        RECT 22.665 2.435 22.915 3.445 ;
  LAYER M1 ;
        RECT 22.665 0.335 22.915 1.345 ;
  LAYER M1 ;
        RECT 23.095 9.575 23.345 13.105 ;
  LAYER M1 ;
        RECT 23.095 3.695 23.345 7.225 ;
  LAYER M1 ;
        RECT 22.235 9.575 22.485 13.105 ;
  LAYER M1 ;
        RECT 22.235 3.695 22.485 7.225 ;
  LAYER M1 ;
        RECT 21.805 9.575 22.055 13.105 ;
  LAYER M1 ;
        RECT 21.805 8.315 22.055 9.325 ;
  LAYER M1 ;
        RECT 21.805 3.695 22.055 7.225 ;
  LAYER M1 ;
        RECT 21.805 2.435 22.055 3.445 ;
  LAYER M1 ;
        RECT 21.805 0.335 22.055 1.345 ;
  LAYER M1 ;
        RECT 21.375 9.575 21.625 13.105 ;
  LAYER M1 ;
        RECT 21.375 3.695 21.625 7.225 ;
  LAYER M1 ;
        RECT 20.945 9.575 21.195 13.105 ;
  LAYER M1 ;
        RECT 20.945 8.315 21.195 9.325 ;
  LAYER M1 ;
        RECT 20.945 3.695 21.195 7.225 ;
  LAYER M1 ;
        RECT 20.945 2.435 21.195 3.445 ;
  LAYER M1 ;
        RECT 20.945 0.335 21.195 1.345 ;
  LAYER M1 ;
        RECT 20.515 9.575 20.765 13.105 ;
  LAYER M1 ;
        RECT 20.515 3.695 20.765 7.225 ;
  LAYER M1 ;
        RECT 20.085 9.575 20.335 13.105 ;
  LAYER M1 ;
        RECT 20.085 8.315 20.335 9.325 ;
  LAYER M1 ;
        RECT 20.085 3.695 20.335 7.225 ;
  LAYER M1 ;
        RECT 20.085 2.435 20.335 3.445 ;
  LAYER M1 ;
        RECT 20.085 0.335 20.335 1.345 ;
  LAYER M1 ;
        RECT 19.655 9.575 19.905 13.105 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M1 ;
        RECT 19.225 9.575 19.475 13.105 ;
  LAYER M1 ;
        RECT 19.225 8.315 19.475 9.325 ;
  LAYER M1 ;
        RECT 19.225 3.695 19.475 7.225 ;
  LAYER M1 ;
        RECT 19.225 2.435 19.475 3.445 ;
  LAYER M1 ;
        RECT 19.225 0.335 19.475 1.345 ;
  LAYER M1 ;
        RECT 18.795 9.575 19.045 13.105 ;
  LAYER M1 ;
        RECT 18.795 3.695 19.045 7.225 ;
  LAYER M1 ;
        RECT 18.365 9.575 18.615 13.105 ;
  LAYER M1 ;
        RECT 18.365 8.315 18.615 9.325 ;
  LAYER M1 ;
        RECT 18.365 3.695 18.615 7.225 ;
  LAYER M1 ;
        RECT 18.365 2.435 18.615 3.445 ;
  LAYER M1 ;
        RECT 18.365 0.335 18.615 1.345 ;
  LAYER M1 ;
        RECT 17.935 9.575 18.185 13.105 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M1 ;
        RECT 17.505 9.575 17.755 13.105 ;
  LAYER M1 ;
        RECT 17.505 8.315 17.755 9.325 ;
  LAYER M1 ;
        RECT 17.505 3.695 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.505 2.435 17.755 3.445 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 1.345 ;
  LAYER M1 ;
        RECT 17.075 9.575 17.325 13.105 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 16.645 9.575 16.895 13.105 ;
  LAYER M1 ;
        RECT 16.645 8.315 16.895 9.325 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 16.215 9.575 16.465 13.105 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 15.785 9.575 16.035 13.105 ;
  LAYER M1 ;
        RECT 15.785 8.315 16.035 9.325 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 15.355 9.575 15.605 13.105 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 14.925 9.575 15.175 13.105 ;
  LAYER M1 ;
        RECT 14.925 8.315 15.175 9.325 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 14.495 9.575 14.745 13.105 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 14.065 9.575 14.315 13.105 ;
  LAYER M1 ;
        RECT 14.065 8.315 14.315 9.325 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 13.635 9.575 13.885 13.105 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 13.205 9.575 13.455 13.105 ;
  LAYER M1 ;
        RECT 13.205 8.315 13.455 9.325 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 9.575 13.025 13.105 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 12.345 9.575 12.595 13.105 ;
  LAYER M1 ;
        RECT 12.345 8.315 12.595 9.325 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 11.915 9.575 12.165 13.105 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 11.485 9.575 11.735 13.105 ;
  LAYER M1 ;
        RECT 11.485 8.315 11.735 9.325 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.055 9.575 11.305 13.105 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 10.625 9.575 10.875 13.105 ;
  LAYER M1 ;
        RECT 10.625 8.315 10.875 9.325 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 10.195 9.575 10.445 13.105 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 9.765 9.575 10.015 13.105 ;
  LAYER M1 ;
        RECT 9.765 8.315 10.015 9.325 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 9.575 9.585 13.105 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 8.905 9.575 9.155 13.105 ;
  LAYER M1 ;
        RECT 8.905 8.315 9.155 9.325 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 8.475 9.575 8.725 13.105 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.045 9.575 8.295 13.105 ;
  LAYER M1 ;
        RECT 8.045 8.315 8.295 9.325 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 7.615 9.575 7.865 13.105 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 7.185 9.575 7.435 13.105 ;
  LAYER M1 ;
        RECT 7.185 8.315 7.435 9.325 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 6.755 9.575 7.005 13.105 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 6.325 9.575 6.575 13.105 ;
  LAYER M1 ;
        RECT 6.325 8.315 6.575 9.325 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 9.575 6.145 13.105 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 5.465 9.575 5.715 13.105 ;
  LAYER M1 ;
        RECT 5.465 8.315 5.715 9.325 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.035 9.575 5.285 13.105 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 4.605 9.575 4.855 13.105 ;
  LAYER M1 ;
        RECT 4.605 8.315 4.855 9.325 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 4.175 9.575 4.425 13.105 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.745 9.575 3.995 13.105 ;
  LAYER M1 ;
        RECT 3.745 8.315 3.995 9.325 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 3.315 9.575 3.565 13.105 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 2.885 9.575 3.135 13.105 ;
  LAYER M1 ;
        RECT 2.885 8.315 3.135 9.325 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 2.455 9.575 2.705 13.105 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.025 9.575 2.275 13.105 ;
  LAYER M1 ;
        RECT 2.025 8.315 2.275 9.325 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 1.595 9.575 1.845 13.105 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 1.165 9.575 1.415 13.105 ;
  LAYER M1 ;
        RECT 1.165 8.315 1.415 9.325 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 9.575 0.985 13.105 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M2 ;
        RECT 1.12 12.88 22.96 13.16 ;
  LAYER M2 ;
        RECT 1.12 8.68 22.96 8.96 ;
  LAYER M2 ;
        RECT 0.69 12.46 23.39 12.74 ;
  LAYER M2 ;
        RECT 1.12 7 22.96 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 22.96 3.08 ;
  LAYER M2 ;
        RECT 0.69 6.58 23.39 6.86 ;
  LAYER M2 ;
        RECT 1.12 0.7 22.96 0.98 ;
  LAYER M3 ;
        RECT 12.33 6.98 12.61 13.18 ;
  LAYER M3 ;
        RECT 11.9 2.78 12.18 8.98 ;
  LAYER M3 ;
        RECT 11.47 0.68 11.75 12.76 ;
  LAYER M1 ;
        RECT 25.245 3.695 25.495 7.225 ;
  LAYER M1 ;
        RECT 25.245 2.435 25.495 3.445 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 1.345 ;
  LAYER M1 ;
        RECT 24.815 3.695 25.065 7.225 ;
  LAYER M1 ;
        RECT 25.675 3.695 25.925 7.225 ;
  LAYER M2 ;
        RECT 24.34 0.7 25.54 0.98 ;
  LAYER M2 ;
        RECT 24.34 7 25.54 7.28 ;
  LAYER M2 ;
        RECT 24.34 2.8 25.54 3.08 ;
  LAYER M2 ;
        RECT 24.77 6.58 25.97 6.86 ;
  LAYER M1 ;
        RECT 27.825 3.695 28.075 7.225 ;
  LAYER M1 ;
        RECT 27.825 2.435 28.075 3.445 ;
  LAYER M1 ;
        RECT 27.825 0.335 28.075 1.345 ;
  LAYER M1 ;
        RECT 28.255 3.695 28.505 7.225 ;
  LAYER M1 ;
        RECT 27.395 3.695 27.645 7.225 ;
  LAYER M2 ;
        RECT 27.78 0.7 28.98 0.98 ;
  LAYER M2 ;
        RECT 27.78 7 28.98 7.28 ;
  LAYER M2 ;
        RECT 27.78 2.8 28.98 3.08 ;
  LAYER M2 ;
        RECT 27.35 6.58 28.55 6.86 ;
  END 
END CURRENT_MIRROR_OTA
