.param w1_2=8.48
.param w3_4=2.5
.param w5_6=67.38
.param w7_8=19.8
.param w9_10=19.00
.param beta=1
.param nf1_2=1
.param nf3_4=1
.param nf5_6=1
.param nf7_8=1
.param nf9_10=1

.param iref_ideal=65u
.param iref_post_layout=65u
