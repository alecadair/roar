MACRO NMOS_S_80601593_X1_Y80
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_80601593_X1_Y80 0 0 ;
  SIZE 2580 BY 472080 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720 260 1000 465100 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 4460 1430 469300 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 471400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 62665 ;
    LAYER M1 ;
      RECT 1165 62915 1415 63925 ;
    LAYER M1 ;
      RECT 1165 65015 1415 68545 ;
    LAYER M1 ;
      RECT 1165 68795 1415 69805 ;
    LAYER M1 ;
      RECT 1165 70895 1415 74425 ;
    LAYER M1 ;
      RECT 1165 74675 1415 75685 ;
    LAYER M1 ;
      RECT 1165 76775 1415 80305 ;
    LAYER M1 ;
      RECT 1165 80555 1415 81565 ;
    LAYER M1 ;
      RECT 1165 82655 1415 86185 ;
    LAYER M1 ;
      RECT 1165 86435 1415 87445 ;
    LAYER M1 ;
      RECT 1165 88535 1415 92065 ;
    LAYER M1 ;
      RECT 1165 92315 1415 93325 ;
    LAYER M1 ;
      RECT 1165 94415 1415 97945 ;
    LAYER M1 ;
      RECT 1165 98195 1415 99205 ;
    LAYER M1 ;
      RECT 1165 100295 1415 103825 ;
    LAYER M1 ;
      RECT 1165 104075 1415 105085 ;
    LAYER M1 ;
      RECT 1165 106175 1415 109705 ;
    LAYER M1 ;
      RECT 1165 109955 1415 110965 ;
    LAYER M1 ;
      RECT 1165 112055 1415 115585 ;
    LAYER M1 ;
      RECT 1165 115835 1415 116845 ;
    LAYER M1 ;
      RECT 1165 117935 1415 121465 ;
    LAYER M1 ;
      RECT 1165 121715 1415 122725 ;
    LAYER M1 ;
      RECT 1165 123815 1415 127345 ;
    LAYER M1 ;
      RECT 1165 127595 1415 128605 ;
    LAYER M1 ;
      RECT 1165 129695 1415 133225 ;
    LAYER M1 ;
      RECT 1165 133475 1415 134485 ;
    LAYER M1 ;
      RECT 1165 135575 1415 139105 ;
    LAYER M1 ;
      RECT 1165 139355 1415 140365 ;
    LAYER M1 ;
      RECT 1165 141455 1415 144985 ;
    LAYER M1 ;
      RECT 1165 145235 1415 146245 ;
    LAYER M1 ;
      RECT 1165 147335 1415 150865 ;
    LAYER M1 ;
      RECT 1165 151115 1415 152125 ;
    LAYER M1 ;
      RECT 1165 153215 1415 156745 ;
    LAYER M1 ;
      RECT 1165 156995 1415 158005 ;
    LAYER M1 ;
      RECT 1165 159095 1415 162625 ;
    LAYER M1 ;
      RECT 1165 162875 1415 163885 ;
    LAYER M1 ;
      RECT 1165 164975 1415 168505 ;
    LAYER M1 ;
      RECT 1165 168755 1415 169765 ;
    LAYER M1 ;
      RECT 1165 170855 1415 174385 ;
    LAYER M1 ;
      RECT 1165 174635 1415 175645 ;
    LAYER M1 ;
      RECT 1165 176735 1415 180265 ;
    LAYER M1 ;
      RECT 1165 180515 1415 181525 ;
    LAYER M1 ;
      RECT 1165 182615 1415 186145 ;
    LAYER M1 ;
      RECT 1165 186395 1415 187405 ;
    LAYER M1 ;
      RECT 1165 188495 1415 192025 ;
    LAYER M1 ;
      RECT 1165 192275 1415 193285 ;
    LAYER M1 ;
      RECT 1165 194375 1415 197905 ;
    LAYER M1 ;
      RECT 1165 198155 1415 199165 ;
    LAYER M1 ;
      RECT 1165 200255 1415 203785 ;
    LAYER M1 ;
      RECT 1165 204035 1415 205045 ;
    LAYER M1 ;
      RECT 1165 206135 1415 209665 ;
    LAYER M1 ;
      RECT 1165 209915 1415 210925 ;
    LAYER M1 ;
      RECT 1165 212015 1415 215545 ;
    LAYER M1 ;
      RECT 1165 215795 1415 216805 ;
    LAYER M1 ;
      RECT 1165 217895 1415 221425 ;
    LAYER M1 ;
      RECT 1165 221675 1415 222685 ;
    LAYER M1 ;
      RECT 1165 223775 1415 227305 ;
    LAYER M1 ;
      RECT 1165 227555 1415 228565 ;
    LAYER M1 ;
      RECT 1165 229655 1415 233185 ;
    LAYER M1 ;
      RECT 1165 233435 1415 234445 ;
    LAYER M1 ;
      RECT 1165 235535 1415 239065 ;
    LAYER M1 ;
      RECT 1165 239315 1415 240325 ;
    LAYER M1 ;
      RECT 1165 241415 1415 244945 ;
    LAYER M1 ;
      RECT 1165 245195 1415 246205 ;
    LAYER M1 ;
      RECT 1165 247295 1415 250825 ;
    LAYER M1 ;
      RECT 1165 251075 1415 252085 ;
    LAYER M1 ;
      RECT 1165 253175 1415 256705 ;
    LAYER M1 ;
      RECT 1165 256955 1415 257965 ;
    LAYER M1 ;
      RECT 1165 259055 1415 262585 ;
    LAYER M1 ;
      RECT 1165 262835 1415 263845 ;
    LAYER M1 ;
      RECT 1165 264935 1415 268465 ;
    LAYER M1 ;
      RECT 1165 268715 1415 269725 ;
    LAYER M1 ;
      RECT 1165 270815 1415 274345 ;
    LAYER M1 ;
      RECT 1165 274595 1415 275605 ;
    LAYER M1 ;
      RECT 1165 276695 1415 280225 ;
    LAYER M1 ;
      RECT 1165 280475 1415 281485 ;
    LAYER M1 ;
      RECT 1165 282575 1415 286105 ;
    LAYER M1 ;
      RECT 1165 286355 1415 287365 ;
    LAYER M1 ;
      RECT 1165 288455 1415 291985 ;
    LAYER M1 ;
      RECT 1165 292235 1415 293245 ;
    LAYER M1 ;
      RECT 1165 294335 1415 297865 ;
    LAYER M1 ;
      RECT 1165 298115 1415 299125 ;
    LAYER M1 ;
      RECT 1165 300215 1415 303745 ;
    LAYER M1 ;
      RECT 1165 303995 1415 305005 ;
    LAYER M1 ;
      RECT 1165 306095 1415 309625 ;
    LAYER M1 ;
      RECT 1165 309875 1415 310885 ;
    LAYER M1 ;
      RECT 1165 311975 1415 315505 ;
    LAYER M1 ;
      RECT 1165 315755 1415 316765 ;
    LAYER M1 ;
      RECT 1165 317855 1415 321385 ;
    LAYER M1 ;
      RECT 1165 321635 1415 322645 ;
    LAYER M1 ;
      RECT 1165 323735 1415 327265 ;
    LAYER M1 ;
      RECT 1165 327515 1415 328525 ;
    LAYER M1 ;
      RECT 1165 329615 1415 333145 ;
    LAYER M1 ;
      RECT 1165 333395 1415 334405 ;
    LAYER M1 ;
      RECT 1165 335495 1415 339025 ;
    LAYER M1 ;
      RECT 1165 339275 1415 340285 ;
    LAYER M1 ;
      RECT 1165 341375 1415 344905 ;
    LAYER M1 ;
      RECT 1165 345155 1415 346165 ;
    LAYER M1 ;
      RECT 1165 347255 1415 350785 ;
    LAYER M1 ;
      RECT 1165 351035 1415 352045 ;
    LAYER M1 ;
      RECT 1165 353135 1415 356665 ;
    LAYER M1 ;
      RECT 1165 356915 1415 357925 ;
    LAYER M1 ;
      RECT 1165 359015 1415 362545 ;
    LAYER M1 ;
      RECT 1165 362795 1415 363805 ;
    LAYER M1 ;
      RECT 1165 364895 1415 368425 ;
    LAYER M1 ;
      RECT 1165 368675 1415 369685 ;
    LAYER M1 ;
      RECT 1165 370775 1415 374305 ;
    LAYER M1 ;
      RECT 1165 374555 1415 375565 ;
    LAYER M1 ;
      RECT 1165 376655 1415 380185 ;
    LAYER M1 ;
      RECT 1165 380435 1415 381445 ;
    LAYER M1 ;
      RECT 1165 382535 1415 386065 ;
    LAYER M1 ;
      RECT 1165 386315 1415 387325 ;
    LAYER M1 ;
      RECT 1165 388415 1415 391945 ;
    LAYER M1 ;
      RECT 1165 392195 1415 393205 ;
    LAYER M1 ;
      RECT 1165 394295 1415 397825 ;
    LAYER M1 ;
      RECT 1165 398075 1415 399085 ;
    LAYER M1 ;
      RECT 1165 400175 1415 403705 ;
    LAYER M1 ;
      RECT 1165 403955 1415 404965 ;
    LAYER M1 ;
      RECT 1165 406055 1415 409585 ;
    LAYER M1 ;
      RECT 1165 409835 1415 410845 ;
    LAYER M1 ;
      RECT 1165 411935 1415 415465 ;
    LAYER M1 ;
      RECT 1165 415715 1415 416725 ;
    LAYER M1 ;
      RECT 1165 417815 1415 421345 ;
    LAYER M1 ;
      RECT 1165 421595 1415 422605 ;
    LAYER M1 ;
      RECT 1165 423695 1415 427225 ;
    LAYER M1 ;
      RECT 1165 427475 1415 428485 ;
    LAYER M1 ;
      RECT 1165 429575 1415 433105 ;
    LAYER M1 ;
      RECT 1165 433355 1415 434365 ;
    LAYER M1 ;
      RECT 1165 435455 1415 438985 ;
    LAYER M1 ;
      RECT 1165 439235 1415 440245 ;
    LAYER M1 ;
      RECT 1165 441335 1415 444865 ;
    LAYER M1 ;
      RECT 1165 445115 1415 446125 ;
    LAYER M1 ;
      RECT 1165 447215 1415 450745 ;
    LAYER M1 ;
      RECT 1165 450995 1415 452005 ;
    LAYER M1 ;
      RECT 1165 453095 1415 456625 ;
    LAYER M1 ;
      RECT 1165 456875 1415 457885 ;
    LAYER M1 ;
      RECT 1165 458975 1415 462505 ;
    LAYER M1 ;
      RECT 1165 462755 1415 463765 ;
    LAYER M1 ;
      RECT 1165 464855 1415 468385 ;
    LAYER M1 ;
      RECT 1165 468635 1415 469645 ;
    LAYER M1 ;
      RECT 1165 470735 1415 471745 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 735 59135 985 62665 ;
    LAYER M1 ;
      RECT 735 65015 985 68545 ;
    LAYER M1 ;
      RECT 735 70895 985 74425 ;
    LAYER M1 ;
      RECT 735 76775 985 80305 ;
    LAYER M1 ;
      RECT 735 82655 985 86185 ;
    LAYER M1 ;
      RECT 735 88535 985 92065 ;
    LAYER M1 ;
      RECT 735 94415 985 97945 ;
    LAYER M1 ;
      RECT 735 100295 985 103825 ;
    LAYER M1 ;
      RECT 735 106175 985 109705 ;
    LAYER M1 ;
      RECT 735 112055 985 115585 ;
    LAYER M1 ;
      RECT 735 117935 985 121465 ;
    LAYER M1 ;
      RECT 735 123815 985 127345 ;
    LAYER M1 ;
      RECT 735 129695 985 133225 ;
    LAYER M1 ;
      RECT 735 135575 985 139105 ;
    LAYER M1 ;
      RECT 735 141455 985 144985 ;
    LAYER M1 ;
      RECT 735 147335 985 150865 ;
    LAYER M1 ;
      RECT 735 153215 985 156745 ;
    LAYER M1 ;
      RECT 735 159095 985 162625 ;
    LAYER M1 ;
      RECT 735 164975 985 168505 ;
    LAYER M1 ;
      RECT 735 170855 985 174385 ;
    LAYER M1 ;
      RECT 735 176735 985 180265 ;
    LAYER M1 ;
      RECT 735 182615 985 186145 ;
    LAYER M1 ;
      RECT 735 188495 985 192025 ;
    LAYER M1 ;
      RECT 735 194375 985 197905 ;
    LAYER M1 ;
      RECT 735 200255 985 203785 ;
    LAYER M1 ;
      RECT 735 206135 985 209665 ;
    LAYER M1 ;
      RECT 735 212015 985 215545 ;
    LAYER M1 ;
      RECT 735 217895 985 221425 ;
    LAYER M1 ;
      RECT 735 223775 985 227305 ;
    LAYER M1 ;
      RECT 735 229655 985 233185 ;
    LAYER M1 ;
      RECT 735 235535 985 239065 ;
    LAYER M1 ;
      RECT 735 241415 985 244945 ;
    LAYER M1 ;
      RECT 735 247295 985 250825 ;
    LAYER M1 ;
      RECT 735 253175 985 256705 ;
    LAYER M1 ;
      RECT 735 259055 985 262585 ;
    LAYER M1 ;
      RECT 735 264935 985 268465 ;
    LAYER M1 ;
      RECT 735 270815 985 274345 ;
    LAYER M1 ;
      RECT 735 276695 985 280225 ;
    LAYER M1 ;
      RECT 735 282575 985 286105 ;
    LAYER M1 ;
      RECT 735 288455 985 291985 ;
    LAYER M1 ;
      RECT 735 294335 985 297865 ;
    LAYER M1 ;
      RECT 735 300215 985 303745 ;
    LAYER M1 ;
      RECT 735 306095 985 309625 ;
    LAYER M1 ;
      RECT 735 311975 985 315505 ;
    LAYER M1 ;
      RECT 735 317855 985 321385 ;
    LAYER M1 ;
      RECT 735 323735 985 327265 ;
    LAYER M1 ;
      RECT 735 329615 985 333145 ;
    LAYER M1 ;
      RECT 735 335495 985 339025 ;
    LAYER M1 ;
      RECT 735 341375 985 344905 ;
    LAYER M1 ;
      RECT 735 347255 985 350785 ;
    LAYER M1 ;
      RECT 735 353135 985 356665 ;
    LAYER M1 ;
      RECT 735 359015 985 362545 ;
    LAYER M1 ;
      RECT 735 364895 985 368425 ;
    LAYER M1 ;
      RECT 735 370775 985 374305 ;
    LAYER M1 ;
      RECT 735 376655 985 380185 ;
    LAYER M1 ;
      RECT 735 382535 985 386065 ;
    LAYER M1 ;
      RECT 735 388415 985 391945 ;
    LAYER M1 ;
      RECT 735 394295 985 397825 ;
    LAYER M1 ;
      RECT 735 400175 985 403705 ;
    LAYER M1 ;
      RECT 735 406055 985 409585 ;
    LAYER M1 ;
      RECT 735 411935 985 415465 ;
    LAYER M1 ;
      RECT 735 417815 985 421345 ;
    LAYER M1 ;
      RECT 735 423695 985 427225 ;
    LAYER M1 ;
      RECT 735 429575 985 433105 ;
    LAYER M1 ;
      RECT 735 435455 985 438985 ;
    LAYER M1 ;
      RECT 735 441335 985 444865 ;
    LAYER M1 ;
      RECT 735 447215 985 450745 ;
    LAYER M1 ;
      RECT 735 453095 985 456625 ;
    LAYER M1 ;
      RECT 735 458975 985 462505 ;
    LAYER M1 ;
      RECT 735 464855 985 468385 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M1 ;
      RECT 1595 59135 1845 62665 ;
    LAYER M1 ;
      RECT 1595 65015 1845 68545 ;
    LAYER M1 ;
      RECT 1595 70895 1845 74425 ;
    LAYER M1 ;
      RECT 1595 76775 1845 80305 ;
    LAYER M1 ;
      RECT 1595 82655 1845 86185 ;
    LAYER M1 ;
      RECT 1595 88535 1845 92065 ;
    LAYER M1 ;
      RECT 1595 94415 1845 97945 ;
    LAYER M1 ;
      RECT 1595 100295 1845 103825 ;
    LAYER M1 ;
      RECT 1595 106175 1845 109705 ;
    LAYER M1 ;
      RECT 1595 112055 1845 115585 ;
    LAYER M1 ;
      RECT 1595 117935 1845 121465 ;
    LAYER M1 ;
      RECT 1595 123815 1845 127345 ;
    LAYER M1 ;
      RECT 1595 129695 1845 133225 ;
    LAYER M1 ;
      RECT 1595 135575 1845 139105 ;
    LAYER M1 ;
      RECT 1595 141455 1845 144985 ;
    LAYER M1 ;
      RECT 1595 147335 1845 150865 ;
    LAYER M1 ;
      RECT 1595 153215 1845 156745 ;
    LAYER M1 ;
      RECT 1595 159095 1845 162625 ;
    LAYER M1 ;
      RECT 1595 164975 1845 168505 ;
    LAYER M1 ;
      RECT 1595 170855 1845 174385 ;
    LAYER M1 ;
      RECT 1595 176735 1845 180265 ;
    LAYER M1 ;
      RECT 1595 182615 1845 186145 ;
    LAYER M1 ;
      RECT 1595 188495 1845 192025 ;
    LAYER M1 ;
      RECT 1595 194375 1845 197905 ;
    LAYER M1 ;
      RECT 1595 200255 1845 203785 ;
    LAYER M1 ;
      RECT 1595 206135 1845 209665 ;
    LAYER M1 ;
      RECT 1595 212015 1845 215545 ;
    LAYER M1 ;
      RECT 1595 217895 1845 221425 ;
    LAYER M1 ;
      RECT 1595 223775 1845 227305 ;
    LAYER M1 ;
      RECT 1595 229655 1845 233185 ;
    LAYER M1 ;
      RECT 1595 235535 1845 239065 ;
    LAYER M1 ;
      RECT 1595 241415 1845 244945 ;
    LAYER M1 ;
      RECT 1595 247295 1845 250825 ;
    LAYER M1 ;
      RECT 1595 253175 1845 256705 ;
    LAYER M1 ;
      RECT 1595 259055 1845 262585 ;
    LAYER M1 ;
      RECT 1595 264935 1845 268465 ;
    LAYER M1 ;
      RECT 1595 270815 1845 274345 ;
    LAYER M1 ;
      RECT 1595 276695 1845 280225 ;
    LAYER M1 ;
      RECT 1595 282575 1845 286105 ;
    LAYER M1 ;
      RECT 1595 288455 1845 291985 ;
    LAYER M1 ;
      RECT 1595 294335 1845 297865 ;
    LAYER M1 ;
      RECT 1595 300215 1845 303745 ;
    LAYER M1 ;
      RECT 1595 306095 1845 309625 ;
    LAYER M1 ;
      RECT 1595 311975 1845 315505 ;
    LAYER M1 ;
      RECT 1595 317855 1845 321385 ;
    LAYER M1 ;
      RECT 1595 323735 1845 327265 ;
    LAYER M1 ;
      RECT 1595 329615 1845 333145 ;
    LAYER M1 ;
      RECT 1595 335495 1845 339025 ;
    LAYER M1 ;
      RECT 1595 341375 1845 344905 ;
    LAYER M1 ;
      RECT 1595 347255 1845 350785 ;
    LAYER M1 ;
      RECT 1595 353135 1845 356665 ;
    LAYER M1 ;
      RECT 1595 359015 1845 362545 ;
    LAYER M1 ;
      RECT 1595 364895 1845 368425 ;
    LAYER M1 ;
      RECT 1595 370775 1845 374305 ;
    LAYER M1 ;
      RECT 1595 376655 1845 380185 ;
    LAYER M1 ;
      RECT 1595 382535 1845 386065 ;
    LAYER M1 ;
      RECT 1595 388415 1845 391945 ;
    LAYER M1 ;
      RECT 1595 394295 1845 397825 ;
    LAYER M1 ;
      RECT 1595 400175 1845 403705 ;
    LAYER M1 ;
      RECT 1595 406055 1845 409585 ;
    LAYER M1 ;
      RECT 1595 411935 1845 415465 ;
    LAYER M1 ;
      RECT 1595 417815 1845 421345 ;
    LAYER M1 ;
      RECT 1595 423695 1845 427225 ;
    LAYER M1 ;
      RECT 1595 429575 1845 433105 ;
    LAYER M1 ;
      RECT 1595 435455 1845 438985 ;
    LAYER M1 ;
      RECT 1595 441335 1845 444865 ;
    LAYER M1 ;
      RECT 1595 447215 1845 450745 ;
    LAYER M1 ;
      RECT 1595 453095 1845 456625 ;
    LAYER M1 ;
      RECT 1595 458975 1845 462505 ;
    LAYER M1 ;
      RECT 1595 464855 1845 468385 ;
    LAYER M2 ;
      RECT 260 280 1460 560 ;
    LAYER M2 ;
      RECT 260 4480 1460 4760 ;
    LAYER M2 ;
      RECT 690 700 1890 980 ;
    LAYER M2 ;
      RECT 260 6160 1460 6440 ;
    LAYER M2 ;
      RECT 260 10360 1460 10640 ;
    LAYER M2 ;
      RECT 690 6580 1890 6860 ;
    LAYER M2 ;
      RECT 260 12040 1460 12320 ;
    LAYER M2 ;
      RECT 260 16240 1460 16520 ;
    LAYER M2 ;
      RECT 690 12460 1890 12740 ;
    LAYER M2 ;
      RECT 260 17920 1460 18200 ;
    LAYER M2 ;
      RECT 260 22120 1460 22400 ;
    LAYER M2 ;
      RECT 690 18340 1890 18620 ;
    LAYER M2 ;
      RECT 260 23800 1460 24080 ;
    LAYER M2 ;
      RECT 260 28000 1460 28280 ;
    LAYER M2 ;
      RECT 690 24220 1890 24500 ;
    LAYER M2 ;
      RECT 260 29680 1460 29960 ;
    LAYER M2 ;
      RECT 260 33880 1460 34160 ;
    LAYER M2 ;
      RECT 690 30100 1890 30380 ;
    LAYER M2 ;
      RECT 260 35560 1460 35840 ;
    LAYER M2 ;
      RECT 260 39760 1460 40040 ;
    LAYER M2 ;
      RECT 690 35980 1890 36260 ;
    LAYER M2 ;
      RECT 260 41440 1460 41720 ;
    LAYER M2 ;
      RECT 260 45640 1460 45920 ;
    LAYER M2 ;
      RECT 690 41860 1890 42140 ;
    LAYER M2 ;
      RECT 260 47320 1460 47600 ;
    LAYER M2 ;
      RECT 260 51520 1460 51800 ;
    LAYER M2 ;
      RECT 690 47740 1890 48020 ;
    LAYER M2 ;
      RECT 260 53200 1460 53480 ;
    LAYER M2 ;
      RECT 260 57400 1460 57680 ;
    LAYER M2 ;
      RECT 690 53620 1890 53900 ;
    LAYER M2 ;
      RECT 260 59080 1460 59360 ;
    LAYER M2 ;
      RECT 260 63280 1460 63560 ;
    LAYER M2 ;
      RECT 690 59500 1890 59780 ;
    LAYER M2 ;
      RECT 260 64960 1460 65240 ;
    LAYER M2 ;
      RECT 260 69160 1460 69440 ;
    LAYER M2 ;
      RECT 690 65380 1890 65660 ;
    LAYER M2 ;
      RECT 260 70840 1460 71120 ;
    LAYER M2 ;
      RECT 260 75040 1460 75320 ;
    LAYER M2 ;
      RECT 690 71260 1890 71540 ;
    LAYER M2 ;
      RECT 260 76720 1460 77000 ;
    LAYER M2 ;
      RECT 260 80920 1460 81200 ;
    LAYER M2 ;
      RECT 690 77140 1890 77420 ;
    LAYER M2 ;
      RECT 260 82600 1460 82880 ;
    LAYER M2 ;
      RECT 260 86800 1460 87080 ;
    LAYER M2 ;
      RECT 690 83020 1890 83300 ;
    LAYER M2 ;
      RECT 260 88480 1460 88760 ;
    LAYER M2 ;
      RECT 260 92680 1460 92960 ;
    LAYER M2 ;
      RECT 690 88900 1890 89180 ;
    LAYER M2 ;
      RECT 260 94360 1460 94640 ;
    LAYER M2 ;
      RECT 260 98560 1460 98840 ;
    LAYER M2 ;
      RECT 690 94780 1890 95060 ;
    LAYER M2 ;
      RECT 260 100240 1460 100520 ;
    LAYER M2 ;
      RECT 260 104440 1460 104720 ;
    LAYER M2 ;
      RECT 690 100660 1890 100940 ;
    LAYER M2 ;
      RECT 260 106120 1460 106400 ;
    LAYER M2 ;
      RECT 260 110320 1460 110600 ;
    LAYER M2 ;
      RECT 690 106540 1890 106820 ;
    LAYER M2 ;
      RECT 260 112000 1460 112280 ;
    LAYER M2 ;
      RECT 260 116200 1460 116480 ;
    LAYER M2 ;
      RECT 690 112420 1890 112700 ;
    LAYER M2 ;
      RECT 260 117880 1460 118160 ;
    LAYER M2 ;
      RECT 260 122080 1460 122360 ;
    LAYER M2 ;
      RECT 690 118300 1890 118580 ;
    LAYER M2 ;
      RECT 260 123760 1460 124040 ;
    LAYER M2 ;
      RECT 260 127960 1460 128240 ;
    LAYER M2 ;
      RECT 690 124180 1890 124460 ;
    LAYER M2 ;
      RECT 260 129640 1460 129920 ;
    LAYER M2 ;
      RECT 260 133840 1460 134120 ;
    LAYER M2 ;
      RECT 690 130060 1890 130340 ;
    LAYER M2 ;
      RECT 260 135520 1460 135800 ;
    LAYER M2 ;
      RECT 260 139720 1460 140000 ;
    LAYER M2 ;
      RECT 690 135940 1890 136220 ;
    LAYER M2 ;
      RECT 260 141400 1460 141680 ;
    LAYER M2 ;
      RECT 260 145600 1460 145880 ;
    LAYER M2 ;
      RECT 690 141820 1890 142100 ;
    LAYER M2 ;
      RECT 260 147280 1460 147560 ;
    LAYER M2 ;
      RECT 260 151480 1460 151760 ;
    LAYER M2 ;
      RECT 690 147700 1890 147980 ;
    LAYER M2 ;
      RECT 260 153160 1460 153440 ;
    LAYER M2 ;
      RECT 260 157360 1460 157640 ;
    LAYER M2 ;
      RECT 690 153580 1890 153860 ;
    LAYER M2 ;
      RECT 260 159040 1460 159320 ;
    LAYER M2 ;
      RECT 260 163240 1460 163520 ;
    LAYER M2 ;
      RECT 690 159460 1890 159740 ;
    LAYER M2 ;
      RECT 260 164920 1460 165200 ;
    LAYER M2 ;
      RECT 260 169120 1460 169400 ;
    LAYER M2 ;
      RECT 690 165340 1890 165620 ;
    LAYER M2 ;
      RECT 260 170800 1460 171080 ;
    LAYER M2 ;
      RECT 260 175000 1460 175280 ;
    LAYER M2 ;
      RECT 690 171220 1890 171500 ;
    LAYER M2 ;
      RECT 260 176680 1460 176960 ;
    LAYER M2 ;
      RECT 260 180880 1460 181160 ;
    LAYER M2 ;
      RECT 690 177100 1890 177380 ;
    LAYER M2 ;
      RECT 260 182560 1460 182840 ;
    LAYER M2 ;
      RECT 260 186760 1460 187040 ;
    LAYER M2 ;
      RECT 690 182980 1890 183260 ;
    LAYER M2 ;
      RECT 260 188440 1460 188720 ;
    LAYER M2 ;
      RECT 260 192640 1460 192920 ;
    LAYER M2 ;
      RECT 690 188860 1890 189140 ;
    LAYER M2 ;
      RECT 260 194320 1460 194600 ;
    LAYER M2 ;
      RECT 260 198520 1460 198800 ;
    LAYER M2 ;
      RECT 690 194740 1890 195020 ;
    LAYER M2 ;
      RECT 260 200200 1460 200480 ;
    LAYER M2 ;
      RECT 260 204400 1460 204680 ;
    LAYER M2 ;
      RECT 690 200620 1890 200900 ;
    LAYER M2 ;
      RECT 260 206080 1460 206360 ;
    LAYER M2 ;
      RECT 260 210280 1460 210560 ;
    LAYER M2 ;
      RECT 690 206500 1890 206780 ;
    LAYER M2 ;
      RECT 260 211960 1460 212240 ;
    LAYER M2 ;
      RECT 260 216160 1460 216440 ;
    LAYER M2 ;
      RECT 690 212380 1890 212660 ;
    LAYER M2 ;
      RECT 260 217840 1460 218120 ;
    LAYER M2 ;
      RECT 260 222040 1460 222320 ;
    LAYER M2 ;
      RECT 690 218260 1890 218540 ;
    LAYER M2 ;
      RECT 260 223720 1460 224000 ;
    LAYER M2 ;
      RECT 260 227920 1460 228200 ;
    LAYER M2 ;
      RECT 690 224140 1890 224420 ;
    LAYER M2 ;
      RECT 260 229600 1460 229880 ;
    LAYER M2 ;
      RECT 260 233800 1460 234080 ;
    LAYER M2 ;
      RECT 690 230020 1890 230300 ;
    LAYER M2 ;
      RECT 260 235480 1460 235760 ;
    LAYER M2 ;
      RECT 260 239680 1460 239960 ;
    LAYER M2 ;
      RECT 690 235900 1890 236180 ;
    LAYER M2 ;
      RECT 260 241360 1460 241640 ;
    LAYER M2 ;
      RECT 260 245560 1460 245840 ;
    LAYER M2 ;
      RECT 690 241780 1890 242060 ;
    LAYER M2 ;
      RECT 260 247240 1460 247520 ;
    LAYER M2 ;
      RECT 260 251440 1460 251720 ;
    LAYER M2 ;
      RECT 690 247660 1890 247940 ;
    LAYER M2 ;
      RECT 260 253120 1460 253400 ;
    LAYER M2 ;
      RECT 260 257320 1460 257600 ;
    LAYER M2 ;
      RECT 690 253540 1890 253820 ;
    LAYER M2 ;
      RECT 260 259000 1460 259280 ;
    LAYER M2 ;
      RECT 260 263200 1460 263480 ;
    LAYER M2 ;
      RECT 690 259420 1890 259700 ;
    LAYER M2 ;
      RECT 260 264880 1460 265160 ;
    LAYER M2 ;
      RECT 260 269080 1460 269360 ;
    LAYER M2 ;
      RECT 690 265300 1890 265580 ;
    LAYER M2 ;
      RECT 260 270760 1460 271040 ;
    LAYER M2 ;
      RECT 260 274960 1460 275240 ;
    LAYER M2 ;
      RECT 690 271180 1890 271460 ;
    LAYER M2 ;
      RECT 260 276640 1460 276920 ;
    LAYER M2 ;
      RECT 260 280840 1460 281120 ;
    LAYER M2 ;
      RECT 690 277060 1890 277340 ;
    LAYER M2 ;
      RECT 260 282520 1460 282800 ;
    LAYER M2 ;
      RECT 260 286720 1460 287000 ;
    LAYER M2 ;
      RECT 690 282940 1890 283220 ;
    LAYER M2 ;
      RECT 260 288400 1460 288680 ;
    LAYER M2 ;
      RECT 260 292600 1460 292880 ;
    LAYER M2 ;
      RECT 690 288820 1890 289100 ;
    LAYER M2 ;
      RECT 260 294280 1460 294560 ;
    LAYER M2 ;
      RECT 260 298480 1460 298760 ;
    LAYER M2 ;
      RECT 690 294700 1890 294980 ;
    LAYER M2 ;
      RECT 260 300160 1460 300440 ;
    LAYER M2 ;
      RECT 260 304360 1460 304640 ;
    LAYER M2 ;
      RECT 690 300580 1890 300860 ;
    LAYER M2 ;
      RECT 260 306040 1460 306320 ;
    LAYER M2 ;
      RECT 260 310240 1460 310520 ;
    LAYER M2 ;
      RECT 690 306460 1890 306740 ;
    LAYER M2 ;
      RECT 260 311920 1460 312200 ;
    LAYER M2 ;
      RECT 260 316120 1460 316400 ;
    LAYER M2 ;
      RECT 690 312340 1890 312620 ;
    LAYER M2 ;
      RECT 260 317800 1460 318080 ;
    LAYER M2 ;
      RECT 260 322000 1460 322280 ;
    LAYER M2 ;
      RECT 690 318220 1890 318500 ;
    LAYER M2 ;
      RECT 260 323680 1460 323960 ;
    LAYER M2 ;
      RECT 260 327880 1460 328160 ;
    LAYER M2 ;
      RECT 690 324100 1890 324380 ;
    LAYER M2 ;
      RECT 260 329560 1460 329840 ;
    LAYER M2 ;
      RECT 260 333760 1460 334040 ;
    LAYER M2 ;
      RECT 690 329980 1890 330260 ;
    LAYER M2 ;
      RECT 260 335440 1460 335720 ;
    LAYER M2 ;
      RECT 260 339640 1460 339920 ;
    LAYER M2 ;
      RECT 690 335860 1890 336140 ;
    LAYER M2 ;
      RECT 260 341320 1460 341600 ;
    LAYER M2 ;
      RECT 260 345520 1460 345800 ;
    LAYER M2 ;
      RECT 690 341740 1890 342020 ;
    LAYER M2 ;
      RECT 260 347200 1460 347480 ;
    LAYER M2 ;
      RECT 260 351400 1460 351680 ;
    LAYER M2 ;
      RECT 690 347620 1890 347900 ;
    LAYER M2 ;
      RECT 260 353080 1460 353360 ;
    LAYER M2 ;
      RECT 260 357280 1460 357560 ;
    LAYER M2 ;
      RECT 690 353500 1890 353780 ;
    LAYER M2 ;
      RECT 260 358960 1460 359240 ;
    LAYER M2 ;
      RECT 260 363160 1460 363440 ;
    LAYER M2 ;
      RECT 690 359380 1890 359660 ;
    LAYER M2 ;
      RECT 260 364840 1460 365120 ;
    LAYER M2 ;
      RECT 260 369040 1460 369320 ;
    LAYER M2 ;
      RECT 690 365260 1890 365540 ;
    LAYER M2 ;
      RECT 260 370720 1460 371000 ;
    LAYER M2 ;
      RECT 260 374920 1460 375200 ;
    LAYER M2 ;
      RECT 690 371140 1890 371420 ;
    LAYER M2 ;
      RECT 260 376600 1460 376880 ;
    LAYER M2 ;
      RECT 260 380800 1460 381080 ;
    LAYER M2 ;
      RECT 690 377020 1890 377300 ;
    LAYER M2 ;
      RECT 260 382480 1460 382760 ;
    LAYER M2 ;
      RECT 260 386680 1460 386960 ;
    LAYER M2 ;
      RECT 690 382900 1890 383180 ;
    LAYER M2 ;
      RECT 260 388360 1460 388640 ;
    LAYER M2 ;
      RECT 260 392560 1460 392840 ;
    LAYER M2 ;
      RECT 690 388780 1890 389060 ;
    LAYER M2 ;
      RECT 260 394240 1460 394520 ;
    LAYER M2 ;
      RECT 260 398440 1460 398720 ;
    LAYER M2 ;
      RECT 690 394660 1890 394940 ;
    LAYER M2 ;
      RECT 260 400120 1460 400400 ;
    LAYER M2 ;
      RECT 260 404320 1460 404600 ;
    LAYER M2 ;
      RECT 690 400540 1890 400820 ;
    LAYER M2 ;
      RECT 260 406000 1460 406280 ;
    LAYER M2 ;
      RECT 260 410200 1460 410480 ;
    LAYER M2 ;
      RECT 690 406420 1890 406700 ;
    LAYER M2 ;
      RECT 260 411880 1460 412160 ;
    LAYER M2 ;
      RECT 260 416080 1460 416360 ;
    LAYER M2 ;
      RECT 690 412300 1890 412580 ;
    LAYER M2 ;
      RECT 260 417760 1460 418040 ;
    LAYER M2 ;
      RECT 260 421960 1460 422240 ;
    LAYER M2 ;
      RECT 690 418180 1890 418460 ;
    LAYER M2 ;
      RECT 260 423640 1460 423920 ;
    LAYER M2 ;
      RECT 260 427840 1460 428120 ;
    LAYER M2 ;
      RECT 690 424060 1890 424340 ;
    LAYER M2 ;
      RECT 260 429520 1460 429800 ;
    LAYER M2 ;
      RECT 260 433720 1460 434000 ;
    LAYER M2 ;
      RECT 690 429940 1890 430220 ;
    LAYER M2 ;
      RECT 260 435400 1460 435680 ;
    LAYER M2 ;
      RECT 260 439600 1460 439880 ;
    LAYER M2 ;
      RECT 690 435820 1890 436100 ;
    LAYER M2 ;
      RECT 260 441280 1460 441560 ;
    LAYER M2 ;
      RECT 260 445480 1460 445760 ;
    LAYER M2 ;
      RECT 690 441700 1890 441980 ;
    LAYER M2 ;
      RECT 260 447160 1460 447440 ;
    LAYER M2 ;
      RECT 260 451360 1460 451640 ;
    LAYER M2 ;
      RECT 690 447580 1890 447860 ;
    LAYER M2 ;
      RECT 260 453040 1460 453320 ;
    LAYER M2 ;
      RECT 260 457240 1460 457520 ;
    LAYER M2 ;
      RECT 690 453460 1890 453740 ;
    LAYER M2 ;
      RECT 260 458920 1460 459200 ;
    LAYER M2 ;
      RECT 260 463120 1460 463400 ;
    LAYER M2 ;
      RECT 690 459340 1890 459620 ;
    LAYER M2 ;
      RECT 260 464800 1460 465080 ;
    LAYER M2 ;
      RECT 260 469000 1460 469280 ;
    LAYER M2 ;
      RECT 690 471100 1890 471380 ;
    LAYER M2 ;
      RECT 690 465220 1890 465500 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53255 1375 53425 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59135 1375 59305 ;
    LAYER V1 ;
      RECT 1205 63335 1375 63505 ;
    LAYER V1 ;
      RECT 1205 65015 1375 65185 ;
    LAYER V1 ;
      RECT 1205 69215 1375 69385 ;
    LAYER V1 ;
      RECT 1205 70895 1375 71065 ;
    LAYER V1 ;
      RECT 1205 75095 1375 75265 ;
    LAYER V1 ;
      RECT 1205 76775 1375 76945 ;
    LAYER V1 ;
      RECT 1205 80975 1375 81145 ;
    LAYER V1 ;
      RECT 1205 82655 1375 82825 ;
    LAYER V1 ;
      RECT 1205 86855 1375 87025 ;
    LAYER V1 ;
      RECT 1205 88535 1375 88705 ;
    LAYER V1 ;
      RECT 1205 92735 1375 92905 ;
    LAYER V1 ;
      RECT 1205 94415 1375 94585 ;
    LAYER V1 ;
      RECT 1205 98615 1375 98785 ;
    LAYER V1 ;
      RECT 1205 100295 1375 100465 ;
    LAYER V1 ;
      RECT 1205 104495 1375 104665 ;
    LAYER V1 ;
      RECT 1205 106175 1375 106345 ;
    LAYER V1 ;
      RECT 1205 110375 1375 110545 ;
    LAYER V1 ;
      RECT 1205 112055 1375 112225 ;
    LAYER V1 ;
      RECT 1205 116255 1375 116425 ;
    LAYER V1 ;
      RECT 1205 117935 1375 118105 ;
    LAYER V1 ;
      RECT 1205 122135 1375 122305 ;
    LAYER V1 ;
      RECT 1205 123815 1375 123985 ;
    LAYER V1 ;
      RECT 1205 128015 1375 128185 ;
    LAYER V1 ;
      RECT 1205 129695 1375 129865 ;
    LAYER V1 ;
      RECT 1205 133895 1375 134065 ;
    LAYER V1 ;
      RECT 1205 135575 1375 135745 ;
    LAYER V1 ;
      RECT 1205 139775 1375 139945 ;
    LAYER V1 ;
      RECT 1205 141455 1375 141625 ;
    LAYER V1 ;
      RECT 1205 145655 1375 145825 ;
    LAYER V1 ;
      RECT 1205 147335 1375 147505 ;
    LAYER V1 ;
      RECT 1205 151535 1375 151705 ;
    LAYER V1 ;
      RECT 1205 153215 1375 153385 ;
    LAYER V1 ;
      RECT 1205 157415 1375 157585 ;
    LAYER V1 ;
      RECT 1205 159095 1375 159265 ;
    LAYER V1 ;
      RECT 1205 163295 1375 163465 ;
    LAYER V1 ;
      RECT 1205 164975 1375 165145 ;
    LAYER V1 ;
      RECT 1205 169175 1375 169345 ;
    LAYER V1 ;
      RECT 1205 170855 1375 171025 ;
    LAYER V1 ;
      RECT 1205 175055 1375 175225 ;
    LAYER V1 ;
      RECT 1205 176735 1375 176905 ;
    LAYER V1 ;
      RECT 1205 180935 1375 181105 ;
    LAYER V1 ;
      RECT 1205 182615 1375 182785 ;
    LAYER V1 ;
      RECT 1205 186815 1375 186985 ;
    LAYER V1 ;
      RECT 1205 188495 1375 188665 ;
    LAYER V1 ;
      RECT 1205 192695 1375 192865 ;
    LAYER V1 ;
      RECT 1205 194375 1375 194545 ;
    LAYER V1 ;
      RECT 1205 198575 1375 198745 ;
    LAYER V1 ;
      RECT 1205 200255 1375 200425 ;
    LAYER V1 ;
      RECT 1205 204455 1375 204625 ;
    LAYER V1 ;
      RECT 1205 206135 1375 206305 ;
    LAYER V1 ;
      RECT 1205 210335 1375 210505 ;
    LAYER V1 ;
      RECT 1205 212015 1375 212185 ;
    LAYER V1 ;
      RECT 1205 216215 1375 216385 ;
    LAYER V1 ;
      RECT 1205 217895 1375 218065 ;
    LAYER V1 ;
      RECT 1205 222095 1375 222265 ;
    LAYER V1 ;
      RECT 1205 223775 1375 223945 ;
    LAYER V1 ;
      RECT 1205 227975 1375 228145 ;
    LAYER V1 ;
      RECT 1205 229655 1375 229825 ;
    LAYER V1 ;
      RECT 1205 233855 1375 234025 ;
    LAYER V1 ;
      RECT 1205 235535 1375 235705 ;
    LAYER V1 ;
      RECT 1205 239735 1375 239905 ;
    LAYER V1 ;
      RECT 1205 241415 1375 241585 ;
    LAYER V1 ;
      RECT 1205 245615 1375 245785 ;
    LAYER V1 ;
      RECT 1205 247295 1375 247465 ;
    LAYER V1 ;
      RECT 1205 251495 1375 251665 ;
    LAYER V1 ;
      RECT 1205 253175 1375 253345 ;
    LAYER V1 ;
      RECT 1205 257375 1375 257545 ;
    LAYER V1 ;
      RECT 1205 259055 1375 259225 ;
    LAYER V1 ;
      RECT 1205 263255 1375 263425 ;
    LAYER V1 ;
      RECT 1205 264935 1375 265105 ;
    LAYER V1 ;
      RECT 1205 269135 1375 269305 ;
    LAYER V1 ;
      RECT 1205 270815 1375 270985 ;
    LAYER V1 ;
      RECT 1205 275015 1375 275185 ;
    LAYER V1 ;
      RECT 1205 276695 1375 276865 ;
    LAYER V1 ;
      RECT 1205 280895 1375 281065 ;
    LAYER V1 ;
      RECT 1205 282575 1375 282745 ;
    LAYER V1 ;
      RECT 1205 286775 1375 286945 ;
    LAYER V1 ;
      RECT 1205 288455 1375 288625 ;
    LAYER V1 ;
      RECT 1205 292655 1375 292825 ;
    LAYER V1 ;
      RECT 1205 294335 1375 294505 ;
    LAYER V1 ;
      RECT 1205 298535 1375 298705 ;
    LAYER V1 ;
      RECT 1205 300215 1375 300385 ;
    LAYER V1 ;
      RECT 1205 304415 1375 304585 ;
    LAYER V1 ;
      RECT 1205 306095 1375 306265 ;
    LAYER V1 ;
      RECT 1205 310295 1375 310465 ;
    LAYER V1 ;
      RECT 1205 311975 1375 312145 ;
    LAYER V1 ;
      RECT 1205 316175 1375 316345 ;
    LAYER V1 ;
      RECT 1205 317855 1375 318025 ;
    LAYER V1 ;
      RECT 1205 322055 1375 322225 ;
    LAYER V1 ;
      RECT 1205 323735 1375 323905 ;
    LAYER V1 ;
      RECT 1205 327935 1375 328105 ;
    LAYER V1 ;
      RECT 1205 329615 1375 329785 ;
    LAYER V1 ;
      RECT 1205 333815 1375 333985 ;
    LAYER V1 ;
      RECT 1205 335495 1375 335665 ;
    LAYER V1 ;
      RECT 1205 339695 1375 339865 ;
    LAYER V1 ;
      RECT 1205 341375 1375 341545 ;
    LAYER V1 ;
      RECT 1205 345575 1375 345745 ;
    LAYER V1 ;
      RECT 1205 347255 1375 347425 ;
    LAYER V1 ;
      RECT 1205 351455 1375 351625 ;
    LAYER V1 ;
      RECT 1205 353135 1375 353305 ;
    LAYER V1 ;
      RECT 1205 357335 1375 357505 ;
    LAYER V1 ;
      RECT 1205 359015 1375 359185 ;
    LAYER V1 ;
      RECT 1205 363215 1375 363385 ;
    LAYER V1 ;
      RECT 1205 364895 1375 365065 ;
    LAYER V1 ;
      RECT 1205 369095 1375 369265 ;
    LAYER V1 ;
      RECT 1205 370775 1375 370945 ;
    LAYER V1 ;
      RECT 1205 374975 1375 375145 ;
    LAYER V1 ;
      RECT 1205 376655 1375 376825 ;
    LAYER V1 ;
      RECT 1205 380855 1375 381025 ;
    LAYER V1 ;
      RECT 1205 382535 1375 382705 ;
    LAYER V1 ;
      RECT 1205 386735 1375 386905 ;
    LAYER V1 ;
      RECT 1205 388415 1375 388585 ;
    LAYER V1 ;
      RECT 1205 392615 1375 392785 ;
    LAYER V1 ;
      RECT 1205 394295 1375 394465 ;
    LAYER V1 ;
      RECT 1205 398495 1375 398665 ;
    LAYER V1 ;
      RECT 1205 400175 1375 400345 ;
    LAYER V1 ;
      RECT 1205 404375 1375 404545 ;
    LAYER V1 ;
      RECT 1205 406055 1375 406225 ;
    LAYER V1 ;
      RECT 1205 410255 1375 410425 ;
    LAYER V1 ;
      RECT 1205 411935 1375 412105 ;
    LAYER V1 ;
      RECT 1205 416135 1375 416305 ;
    LAYER V1 ;
      RECT 1205 417815 1375 417985 ;
    LAYER V1 ;
      RECT 1205 422015 1375 422185 ;
    LAYER V1 ;
      RECT 1205 423695 1375 423865 ;
    LAYER V1 ;
      RECT 1205 427895 1375 428065 ;
    LAYER V1 ;
      RECT 1205 429575 1375 429745 ;
    LAYER V1 ;
      RECT 1205 433775 1375 433945 ;
    LAYER V1 ;
      RECT 1205 435455 1375 435625 ;
    LAYER V1 ;
      RECT 1205 439655 1375 439825 ;
    LAYER V1 ;
      RECT 1205 441335 1375 441505 ;
    LAYER V1 ;
      RECT 1205 445535 1375 445705 ;
    LAYER V1 ;
      RECT 1205 447215 1375 447385 ;
    LAYER V1 ;
      RECT 1205 451415 1375 451585 ;
    LAYER V1 ;
      RECT 1205 453095 1375 453265 ;
    LAYER V1 ;
      RECT 1205 457295 1375 457465 ;
    LAYER V1 ;
      RECT 1205 458975 1375 459145 ;
    LAYER V1 ;
      RECT 1205 463175 1375 463345 ;
    LAYER V1 ;
      RECT 1205 464855 1375 465025 ;
    LAYER V1 ;
      RECT 1205 469055 1375 469225 ;
    LAYER V1 ;
      RECT 1205 471155 1375 471325 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 775 53675 945 53845 ;
    LAYER V1 ;
      RECT 775 59555 945 59725 ;
    LAYER V1 ;
      RECT 775 65435 945 65605 ;
    LAYER V1 ;
      RECT 775 71315 945 71485 ;
    LAYER V1 ;
      RECT 775 77195 945 77365 ;
    LAYER V1 ;
      RECT 775 83075 945 83245 ;
    LAYER V1 ;
      RECT 775 88955 945 89125 ;
    LAYER V1 ;
      RECT 775 94835 945 95005 ;
    LAYER V1 ;
      RECT 775 100715 945 100885 ;
    LAYER V1 ;
      RECT 775 106595 945 106765 ;
    LAYER V1 ;
      RECT 775 112475 945 112645 ;
    LAYER V1 ;
      RECT 775 118355 945 118525 ;
    LAYER V1 ;
      RECT 775 124235 945 124405 ;
    LAYER V1 ;
      RECT 775 130115 945 130285 ;
    LAYER V1 ;
      RECT 775 135995 945 136165 ;
    LAYER V1 ;
      RECT 775 141875 945 142045 ;
    LAYER V1 ;
      RECT 775 147755 945 147925 ;
    LAYER V1 ;
      RECT 775 153635 945 153805 ;
    LAYER V1 ;
      RECT 775 159515 945 159685 ;
    LAYER V1 ;
      RECT 775 165395 945 165565 ;
    LAYER V1 ;
      RECT 775 171275 945 171445 ;
    LAYER V1 ;
      RECT 775 177155 945 177325 ;
    LAYER V1 ;
      RECT 775 183035 945 183205 ;
    LAYER V1 ;
      RECT 775 188915 945 189085 ;
    LAYER V1 ;
      RECT 775 194795 945 194965 ;
    LAYER V1 ;
      RECT 775 200675 945 200845 ;
    LAYER V1 ;
      RECT 775 206555 945 206725 ;
    LAYER V1 ;
      RECT 775 212435 945 212605 ;
    LAYER V1 ;
      RECT 775 218315 945 218485 ;
    LAYER V1 ;
      RECT 775 224195 945 224365 ;
    LAYER V1 ;
      RECT 775 230075 945 230245 ;
    LAYER V1 ;
      RECT 775 235955 945 236125 ;
    LAYER V1 ;
      RECT 775 241835 945 242005 ;
    LAYER V1 ;
      RECT 775 247715 945 247885 ;
    LAYER V1 ;
      RECT 775 253595 945 253765 ;
    LAYER V1 ;
      RECT 775 259475 945 259645 ;
    LAYER V1 ;
      RECT 775 265355 945 265525 ;
    LAYER V1 ;
      RECT 775 271235 945 271405 ;
    LAYER V1 ;
      RECT 775 277115 945 277285 ;
    LAYER V1 ;
      RECT 775 282995 945 283165 ;
    LAYER V1 ;
      RECT 775 288875 945 289045 ;
    LAYER V1 ;
      RECT 775 294755 945 294925 ;
    LAYER V1 ;
      RECT 775 300635 945 300805 ;
    LAYER V1 ;
      RECT 775 306515 945 306685 ;
    LAYER V1 ;
      RECT 775 312395 945 312565 ;
    LAYER V1 ;
      RECT 775 318275 945 318445 ;
    LAYER V1 ;
      RECT 775 324155 945 324325 ;
    LAYER V1 ;
      RECT 775 330035 945 330205 ;
    LAYER V1 ;
      RECT 775 335915 945 336085 ;
    LAYER V1 ;
      RECT 775 341795 945 341965 ;
    LAYER V1 ;
      RECT 775 347675 945 347845 ;
    LAYER V1 ;
      RECT 775 353555 945 353725 ;
    LAYER V1 ;
      RECT 775 359435 945 359605 ;
    LAYER V1 ;
      RECT 775 365315 945 365485 ;
    LAYER V1 ;
      RECT 775 371195 945 371365 ;
    LAYER V1 ;
      RECT 775 377075 945 377245 ;
    LAYER V1 ;
      RECT 775 382955 945 383125 ;
    LAYER V1 ;
      RECT 775 388835 945 389005 ;
    LAYER V1 ;
      RECT 775 394715 945 394885 ;
    LAYER V1 ;
      RECT 775 400595 945 400765 ;
    LAYER V1 ;
      RECT 775 406475 945 406645 ;
    LAYER V1 ;
      RECT 775 412355 945 412525 ;
    LAYER V1 ;
      RECT 775 418235 945 418405 ;
    LAYER V1 ;
      RECT 775 424115 945 424285 ;
    LAYER V1 ;
      RECT 775 429995 945 430165 ;
    LAYER V1 ;
      RECT 775 435875 945 436045 ;
    LAYER V1 ;
      RECT 775 441755 945 441925 ;
    LAYER V1 ;
      RECT 775 447635 945 447805 ;
    LAYER V1 ;
      RECT 775 453515 945 453685 ;
    LAYER V1 ;
      RECT 775 459395 945 459565 ;
    LAYER V1 ;
      RECT 775 465275 945 465445 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 1635 53675 1805 53845 ;
    LAYER V1 ;
      RECT 1635 59555 1805 59725 ;
    LAYER V1 ;
      RECT 1635 65435 1805 65605 ;
    LAYER V1 ;
      RECT 1635 71315 1805 71485 ;
    LAYER V1 ;
      RECT 1635 77195 1805 77365 ;
    LAYER V1 ;
      RECT 1635 83075 1805 83245 ;
    LAYER V1 ;
      RECT 1635 88955 1805 89125 ;
    LAYER V1 ;
      RECT 1635 94835 1805 95005 ;
    LAYER V1 ;
      RECT 1635 100715 1805 100885 ;
    LAYER V1 ;
      RECT 1635 106595 1805 106765 ;
    LAYER V1 ;
      RECT 1635 112475 1805 112645 ;
    LAYER V1 ;
      RECT 1635 118355 1805 118525 ;
    LAYER V1 ;
      RECT 1635 124235 1805 124405 ;
    LAYER V1 ;
      RECT 1635 130115 1805 130285 ;
    LAYER V1 ;
      RECT 1635 135995 1805 136165 ;
    LAYER V1 ;
      RECT 1635 141875 1805 142045 ;
    LAYER V1 ;
      RECT 1635 147755 1805 147925 ;
    LAYER V1 ;
      RECT 1635 153635 1805 153805 ;
    LAYER V1 ;
      RECT 1635 159515 1805 159685 ;
    LAYER V1 ;
      RECT 1635 165395 1805 165565 ;
    LAYER V1 ;
      RECT 1635 171275 1805 171445 ;
    LAYER V1 ;
      RECT 1635 177155 1805 177325 ;
    LAYER V1 ;
      RECT 1635 183035 1805 183205 ;
    LAYER V1 ;
      RECT 1635 188915 1805 189085 ;
    LAYER V1 ;
      RECT 1635 194795 1805 194965 ;
    LAYER V1 ;
      RECT 1635 200675 1805 200845 ;
    LAYER V1 ;
      RECT 1635 206555 1805 206725 ;
    LAYER V1 ;
      RECT 1635 212435 1805 212605 ;
    LAYER V1 ;
      RECT 1635 218315 1805 218485 ;
    LAYER V1 ;
      RECT 1635 224195 1805 224365 ;
    LAYER V1 ;
      RECT 1635 230075 1805 230245 ;
    LAYER V1 ;
      RECT 1635 235955 1805 236125 ;
    LAYER V1 ;
      RECT 1635 241835 1805 242005 ;
    LAYER V1 ;
      RECT 1635 247715 1805 247885 ;
    LAYER V1 ;
      RECT 1635 253595 1805 253765 ;
    LAYER V1 ;
      RECT 1635 259475 1805 259645 ;
    LAYER V1 ;
      RECT 1635 265355 1805 265525 ;
    LAYER V1 ;
      RECT 1635 271235 1805 271405 ;
    LAYER V1 ;
      RECT 1635 277115 1805 277285 ;
    LAYER V1 ;
      RECT 1635 282995 1805 283165 ;
    LAYER V1 ;
      RECT 1635 288875 1805 289045 ;
    LAYER V1 ;
      RECT 1635 294755 1805 294925 ;
    LAYER V1 ;
      RECT 1635 300635 1805 300805 ;
    LAYER V1 ;
      RECT 1635 306515 1805 306685 ;
    LAYER V1 ;
      RECT 1635 312395 1805 312565 ;
    LAYER V1 ;
      RECT 1635 318275 1805 318445 ;
    LAYER V1 ;
      RECT 1635 324155 1805 324325 ;
    LAYER V1 ;
      RECT 1635 330035 1805 330205 ;
    LAYER V1 ;
      RECT 1635 335915 1805 336085 ;
    LAYER V1 ;
      RECT 1635 341795 1805 341965 ;
    LAYER V1 ;
      RECT 1635 347675 1805 347845 ;
    LAYER V1 ;
      RECT 1635 353555 1805 353725 ;
    LAYER V1 ;
      RECT 1635 359435 1805 359605 ;
    LAYER V1 ;
      RECT 1635 365315 1805 365485 ;
    LAYER V1 ;
      RECT 1635 371195 1805 371365 ;
    LAYER V1 ;
      RECT 1635 377075 1805 377245 ;
    LAYER V1 ;
      RECT 1635 382955 1805 383125 ;
    LAYER V1 ;
      RECT 1635 388835 1805 389005 ;
    LAYER V1 ;
      RECT 1635 394715 1805 394885 ;
    LAYER V1 ;
      RECT 1635 400595 1805 400765 ;
    LAYER V1 ;
      RECT 1635 406475 1805 406645 ;
    LAYER V1 ;
      RECT 1635 412355 1805 412525 ;
    LAYER V1 ;
      RECT 1635 418235 1805 418405 ;
    LAYER V1 ;
      RECT 1635 424115 1805 424285 ;
    LAYER V1 ;
      RECT 1635 429995 1805 430165 ;
    LAYER V1 ;
      RECT 1635 435875 1805 436045 ;
    LAYER V1 ;
      RECT 1635 441755 1805 441925 ;
    LAYER V1 ;
      RECT 1635 447635 1805 447805 ;
    LAYER V1 ;
      RECT 1635 453515 1805 453685 ;
    LAYER V1 ;
      RECT 1635 459395 1805 459565 ;
    LAYER V1 ;
      RECT 1635 465275 1805 465445 ;
    LAYER V2 ;
      RECT 785 345 935 495 ;
    LAYER V2 ;
      RECT 785 6225 935 6375 ;
    LAYER V2 ;
      RECT 785 12105 935 12255 ;
    LAYER V2 ;
      RECT 785 17985 935 18135 ;
    LAYER V2 ;
      RECT 785 23865 935 24015 ;
    LAYER V2 ;
      RECT 785 29745 935 29895 ;
    LAYER V2 ;
      RECT 785 35625 935 35775 ;
    LAYER V2 ;
      RECT 785 41505 935 41655 ;
    LAYER V2 ;
      RECT 785 47385 935 47535 ;
    LAYER V2 ;
      RECT 785 53265 935 53415 ;
    LAYER V2 ;
      RECT 785 59145 935 59295 ;
    LAYER V2 ;
      RECT 785 65025 935 65175 ;
    LAYER V2 ;
      RECT 785 70905 935 71055 ;
    LAYER V2 ;
      RECT 785 76785 935 76935 ;
    LAYER V2 ;
      RECT 785 82665 935 82815 ;
    LAYER V2 ;
      RECT 785 88545 935 88695 ;
    LAYER V2 ;
      RECT 785 94425 935 94575 ;
    LAYER V2 ;
      RECT 785 100305 935 100455 ;
    LAYER V2 ;
      RECT 785 106185 935 106335 ;
    LAYER V2 ;
      RECT 785 112065 935 112215 ;
    LAYER V2 ;
      RECT 785 117945 935 118095 ;
    LAYER V2 ;
      RECT 785 123825 935 123975 ;
    LAYER V2 ;
      RECT 785 129705 935 129855 ;
    LAYER V2 ;
      RECT 785 135585 935 135735 ;
    LAYER V2 ;
      RECT 785 141465 935 141615 ;
    LAYER V2 ;
      RECT 785 147345 935 147495 ;
    LAYER V2 ;
      RECT 785 153225 935 153375 ;
    LAYER V2 ;
      RECT 785 159105 935 159255 ;
    LAYER V2 ;
      RECT 785 164985 935 165135 ;
    LAYER V2 ;
      RECT 785 170865 935 171015 ;
    LAYER V2 ;
      RECT 785 176745 935 176895 ;
    LAYER V2 ;
      RECT 785 182625 935 182775 ;
    LAYER V2 ;
      RECT 785 188505 935 188655 ;
    LAYER V2 ;
      RECT 785 194385 935 194535 ;
    LAYER V2 ;
      RECT 785 200265 935 200415 ;
    LAYER V2 ;
      RECT 785 206145 935 206295 ;
    LAYER V2 ;
      RECT 785 212025 935 212175 ;
    LAYER V2 ;
      RECT 785 217905 935 218055 ;
    LAYER V2 ;
      RECT 785 223785 935 223935 ;
    LAYER V2 ;
      RECT 785 229665 935 229815 ;
    LAYER V2 ;
      RECT 785 235545 935 235695 ;
    LAYER V2 ;
      RECT 785 241425 935 241575 ;
    LAYER V2 ;
      RECT 785 247305 935 247455 ;
    LAYER V2 ;
      RECT 785 253185 935 253335 ;
    LAYER V2 ;
      RECT 785 259065 935 259215 ;
    LAYER V2 ;
      RECT 785 264945 935 265095 ;
    LAYER V2 ;
      RECT 785 270825 935 270975 ;
    LAYER V2 ;
      RECT 785 276705 935 276855 ;
    LAYER V2 ;
      RECT 785 282585 935 282735 ;
    LAYER V2 ;
      RECT 785 288465 935 288615 ;
    LAYER V2 ;
      RECT 785 294345 935 294495 ;
    LAYER V2 ;
      RECT 785 300225 935 300375 ;
    LAYER V2 ;
      RECT 785 306105 935 306255 ;
    LAYER V2 ;
      RECT 785 311985 935 312135 ;
    LAYER V2 ;
      RECT 785 317865 935 318015 ;
    LAYER V2 ;
      RECT 785 323745 935 323895 ;
    LAYER V2 ;
      RECT 785 329625 935 329775 ;
    LAYER V2 ;
      RECT 785 335505 935 335655 ;
    LAYER V2 ;
      RECT 785 341385 935 341535 ;
    LAYER V2 ;
      RECT 785 347265 935 347415 ;
    LAYER V2 ;
      RECT 785 353145 935 353295 ;
    LAYER V2 ;
      RECT 785 359025 935 359175 ;
    LAYER V2 ;
      RECT 785 364905 935 365055 ;
    LAYER V2 ;
      RECT 785 370785 935 370935 ;
    LAYER V2 ;
      RECT 785 376665 935 376815 ;
    LAYER V2 ;
      RECT 785 382545 935 382695 ;
    LAYER V2 ;
      RECT 785 388425 935 388575 ;
    LAYER V2 ;
      RECT 785 394305 935 394455 ;
    LAYER V2 ;
      RECT 785 400185 935 400335 ;
    LAYER V2 ;
      RECT 785 406065 935 406215 ;
    LAYER V2 ;
      RECT 785 411945 935 412095 ;
    LAYER V2 ;
      RECT 785 417825 935 417975 ;
    LAYER V2 ;
      RECT 785 423705 935 423855 ;
    LAYER V2 ;
      RECT 785 429585 935 429735 ;
    LAYER V2 ;
      RECT 785 435465 935 435615 ;
    LAYER V2 ;
      RECT 785 441345 935 441495 ;
    LAYER V2 ;
      RECT 785 447225 935 447375 ;
    LAYER V2 ;
      RECT 785 453105 935 453255 ;
    LAYER V2 ;
      RECT 785 458985 935 459135 ;
    LAYER V2 ;
      RECT 785 464865 935 465015 ;
    LAYER V2 ;
      RECT 1215 4545 1365 4695 ;
    LAYER V2 ;
      RECT 1215 10425 1365 10575 ;
    LAYER V2 ;
      RECT 1215 16305 1365 16455 ;
    LAYER V2 ;
      RECT 1215 22185 1365 22335 ;
    LAYER V2 ;
      RECT 1215 28065 1365 28215 ;
    LAYER V2 ;
      RECT 1215 33945 1365 34095 ;
    LAYER V2 ;
      RECT 1215 39825 1365 39975 ;
    LAYER V2 ;
      RECT 1215 45705 1365 45855 ;
    LAYER V2 ;
      RECT 1215 51585 1365 51735 ;
    LAYER V2 ;
      RECT 1215 57465 1365 57615 ;
    LAYER V2 ;
      RECT 1215 63345 1365 63495 ;
    LAYER V2 ;
      RECT 1215 69225 1365 69375 ;
    LAYER V2 ;
      RECT 1215 75105 1365 75255 ;
    LAYER V2 ;
      RECT 1215 80985 1365 81135 ;
    LAYER V2 ;
      RECT 1215 86865 1365 87015 ;
    LAYER V2 ;
      RECT 1215 92745 1365 92895 ;
    LAYER V2 ;
      RECT 1215 98625 1365 98775 ;
    LAYER V2 ;
      RECT 1215 104505 1365 104655 ;
    LAYER V2 ;
      RECT 1215 110385 1365 110535 ;
    LAYER V2 ;
      RECT 1215 116265 1365 116415 ;
    LAYER V2 ;
      RECT 1215 122145 1365 122295 ;
    LAYER V2 ;
      RECT 1215 128025 1365 128175 ;
    LAYER V2 ;
      RECT 1215 133905 1365 134055 ;
    LAYER V2 ;
      RECT 1215 139785 1365 139935 ;
    LAYER V2 ;
      RECT 1215 145665 1365 145815 ;
    LAYER V2 ;
      RECT 1215 151545 1365 151695 ;
    LAYER V2 ;
      RECT 1215 157425 1365 157575 ;
    LAYER V2 ;
      RECT 1215 163305 1365 163455 ;
    LAYER V2 ;
      RECT 1215 169185 1365 169335 ;
    LAYER V2 ;
      RECT 1215 175065 1365 175215 ;
    LAYER V2 ;
      RECT 1215 180945 1365 181095 ;
    LAYER V2 ;
      RECT 1215 186825 1365 186975 ;
    LAYER V2 ;
      RECT 1215 192705 1365 192855 ;
    LAYER V2 ;
      RECT 1215 198585 1365 198735 ;
    LAYER V2 ;
      RECT 1215 204465 1365 204615 ;
    LAYER V2 ;
      RECT 1215 210345 1365 210495 ;
    LAYER V2 ;
      RECT 1215 216225 1365 216375 ;
    LAYER V2 ;
      RECT 1215 222105 1365 222255 ;
    LAYER V2 ;
      RECT 1215 227985 1365 228135 ;
    LAYER V2 ;
      RECT 1215 233865 1365 234015 ;
    LAYER V2 ;
      RECT 1215 239745 1365 239895 ;
    LAYER V2 ;
      RECT 1215 245625 1365 245775 ;
    LAYER V2 ;
      RECT 1215 251505 1365 251655 ;
    LAYER V2 ;
      RECT 1215 257385 1365 257535 ;
    LAYER V2 ;
      RECT 1215 263265 1365 263415 ;
    LAYER V2 ;
      RECT 1215 269145 1365 269295 ;
    LAYER V2 ;
      RECT 1215 275025 1365 275175 ;
    LAYER V2 ;
      RECT 1215 280905 1365 281055 ;
    LAYER V2 ;
      RECT 1215 286785 1365 286935 ;
    LAYER V2 ;
      RECT 1215 292665 1365 292815 ;
    LAYER V2 ;
      RECT 1215 298545 1365 298695 ;
    LAYER V2 ;
      RECT 1215 304425 1365 304575 ;
    LAYER V2 ;
      RECT 1215 310305 1365 310455 ;
    LAYER V2 ;
      RECT 1215 316185 1365 316335 ;
    LAYER V2 ;
      RECT 1215 322065 1365 322215 ;
    LAYER V2 ;
      RECT 1215 327945 1365 328095 ;
    LAYER V2 ;
      RECT 1215 333825 1365 333975 ;
    LAYER V2 ;
      RECT 1215 339705 1365 339855 ;
    LAYER V2 ;
      RECT 1215 345585 1365 345735 ;
    LAYER V2 ;
      RECT 1215 351465 1365 351615 ;
    LAYER V2 ;
      RECT 1215 357345 1365 357495 ;
    LAYER V2 ;
      RECT 1215 363225 1365 363375 ;
    LAYER V2 ;
      RECT 1215 369105 1365 369255 ;
    LAYER V2 ;
      RECT 1215 374985 1365 375135 ;
    LAYER V2 ;
      RECT 1215 380865 1365 381015 ;
    LAYER V2 ;
      RECT 1215 386745 1365 386895 ;
    LAYER V2 ;
      RECT 1215 392625 1365 392775 ;
    LAYER V2 ;
      RECT 1215 398505 1365 398655 ;
    LAYER V2 ;
      RECT 1215 404385 1365 404535 ;
    LAYER V2 ;
      RECT 1215 410265 1365 410415 ;
    LAYER V2 ;
      RECT 1215 416145 1365 416295 ;
    LAYER V2 ;
      RECT 1215 422025 1365 422175 ;
    LAYER V2 ;
      RECT 1215 427905 1365 428055 ;
    LAYER V2 ;
      RECT 1215 433785 1365 433935 ;
    LAYER V2 ;
      RECT 1215 439665 1365 439815 ;
    LAYER V2 ;
      RECT 1215 445545 1365 445695 ;
    LAYER V2 ;
      RECT 1215 451425 1365 451575 ;
    LAYER V2 ;
      RECT 1215 457305 1365 457455 ;
    LAYER V2 ;
      RECT 1215 463185 1365 463335 ;
    LAYER V2 ;
      RECT 1215 469065 1365 469215 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 6645 1795 6795 ;
    LAYER V2 ;
      RECT 1645 12525 1795 12675 ;
    LAYER V2 ;
      RECT 1645 18405 1795 18555 ;
    LAYER V2 ;
      RECT 1645 24285 1795 24435 ;
    LAYER V2 ;
      RECT 1645 30165 1795 30315 ;
    LAYER V2 ;
      RECT 1645 36045 1795 36195 ;
    LAYER V2 ;
      RECT 1645 41925 1795 42075 ;
    LAYER V2 ;
      RECT 1645 47805 1795 47955 ;
    LAYER V2 ;
      RECT 1645 53685 1795 53835 ;
    LAYER V2 ;
      RECT 1645 59565 1795 59715 ;
    LAYER V2 ;
      RECT 1645 65445 1795 65595 ;
    LAYER V2 ;
      RECT 1645 71325 1795 71475 ;
    LAYER V2 ;
      RECT 1645 77205 1795 77355 ;
    LAYER V2 ;
      RECT 1645 83085 1795 83235 ;
    LAYER V2 ;
      RECT 1645 88965 1795 89115 ;
    LAYER V2 ;
      RECT 1645 94845 1795 94995 ;
    LAYER V2 ;
      RECT 1645 100725 1795 100875 ;
    LAYER V2 ;
      RECT 1645 106605 1795 106755 ;
    LAYER V2 ;
      RECT 1645 112485 1795 112635 ;
    LAYER V2 ;
      RECT 1645 118365 1795 118515 ;
    LAYER V2 ;
      RECT 1645 124245 1795 124395 ;
    LAYER V2 ;
      RECT 1645 130125 1795 130275 ;
    LAYER V2 ;
      RECT 1645 136005 1795 136155 ;
    LAYER V2 ;
      RECT 1645 141885 1795 142035 ;
    LAYER V2 ;
      RECT 1645 147765 1795 147915 ;
    LAYER V2 ;
      RECT 1645 153645 1795 153795 ;
    LAYER V2 ;
      RECT 1645 159525 1795 159675 ;
    LAYER V2 ;
      RECT 1645 165405 1795 165555 ;
    LAYER V2 ;
      RECT 1645 171285 1795 171435 ;
    LAYER V2 ;
      RECT 1645 177165 1795 177315 ;
    LAYER V2 ;
      RECT 1645 183045 1795 183195 ;
    LAYER V2 ;
      RECT 1645 188925 1795 189075 ;
    LAYER V2 ;
      RECT 1645 194805 1795 194955 ;
    LAYER V2 ;
      RECT 1645 200685 1795 200835 ;
    LAYER V2 ;
      RECT 1645 206565 1795 206715 ;
    LAYER V2 ;
      RECT 1645 212445 1795 212595 ;
    LAYER V2 ;
      RECT 1645 218325 1795 218475 ;
    LAYER V2 ;
      RECT 1645 224205 1795 224355 ;
    LAYER V2 ;
      RECT 1645 230085 1795 230235 ;
    LAYER V2 ;
      RECT 1645 235965 1795 236115 ;
    LAYER V2 ;
      RECT 1645 241845 1795 241995 ;
    LAYER V2 ;
      RECT 1645 247725 1795 247875 ;
    LAYER V2 ;
      RECT 1645 253605 1795 253755 ;
    LAYER V2 ;
      RECT 1645 259485 1795 259635 ;
    LAYER V2 ;
      RECT 1645 265365 1795 265515 ;
    LAYER V2 ;
      RECT 1645 271245 1795 271395 ;
    LAYER V2 ;
      RECT 1645 277125 1795 277275 ;
    LAYER V2 ;
      RECT 1645 283005 1795 283155 ;
    LAYER V2 ;
      RECT 1645 288885 1795 289035 ;
    LAYER V2 ;
      RECT 1645 294765 1795 294915 ;
    LAYER V2 ;
      RECT 1645 300645 1795 300795 ;
    LAYER V2 ;
      RECT 1645 306525 1795 306675 ;
    LAYER V2 ;
      RECT 1645 312405 1795 312555 ;
    LAYER V2 ;
      RECT 1645 318285 1795 318435 ;
    LAYER V2 ;
      RECT 1645 324165 1795 324315 ;
    LAYER V2 ;
      RECT 1645 330045 1795 330195 ;
    LAYER V2 ;
      RECT 1645 335925 1795 336075 ;
    LAYER V2 ;
      RECT 1645 341805 1795 341955 ;
    LAYER V2 ;
      RECT 1645 347685 1795 347835 ;
    LAYER V2 ;
      RECT 1645 353565 1795 353715 ;
    LAYER V2 ;
      RECT 1645 359445 1795 359595 ;
    LAYER V2 ;
      RECT 1645 365325 1795 365475 ;
    LAYER V2 ;
      RECT 1645 371205 1795 371355 ;
    LAYER V2 ;
      RECT 1645 377085 1795 377235 ;
    LAYER V2 ;
      RECT 1645 382965 1795 383115 ;
    LAYER V2 ;
      RECT 1645 388845 1795 388995 ;
    LAYER V2 ;
      RECT 1645 394725 1795 394875 ;
    LAYER V2 ;
      RECT 1645 400605 1795 400755 ;
    LAYER V2 ;
      RECT 1645 406485 1795 406635 ;
    LAYER V2 ;
      RECT 1645 412365 1795 412515 ;
    LAYER V2 ;
      RECT 1645 418245 1795 418395 ;
    LAYER V2 ;
      RECT 1645 424125 1795 424275 ;
    LAYER V2 ;
      RECT 1645 430005 1795 430155 ;
    LAYER V2 ;
      RECT 1645 435885 1795 436035 ;
    LAYER V2 ;
      RECT 1645 441765 1795 441915 ;
    LAYER V2 ;
      RECT 1645 447645 1795 447795 ;
    LAYER V2 ;
      RECT 1645 453525 1795 453675 ;
    LAYER V2 ;
      RECT 1645 459405 1795 459555 ;
    LAYER V2 ;
      RECT 1645 465285 1795 465435 ;
    LAYER V2 ;
      RECT 1645 471165 1795 471315 ;
  END
END NMOS_S_80601593_X1_Y80
