MACRO NMOS_S_80601593_X8_Y10
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_80601593_X8_Y10 0 0 ;
  SIZE 8600 BY 60480 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3730 260 4010 53500 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 4160 4460 4440 57700 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 4590 680 4870 59800 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 60145 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 33265 ;
    LAYER M1 ;
      RECT 2025 33515 2275 34525 ;
    LAYER M1 ;
      RECT 2025 35615 2275 39145 ;
    LAYER M1 ;
      RECT 2025 39395 2275 40405 ;
    LAYER M1 ;
      RECT 2025 41495 2275 45025 ;
    LAYER M1 ;
      RECT 2025 45275 2275 46285 ;
    LAYER M1 ;
      RECT 2025 47375 2275 50905 ;
    LAYER M1 ;
      RECT 2025 51155 2275 52165 ;
    LAYER M1 ;
      RECT 2025 53255 2275 56785 ;
    LAYER M1 ;
      RECT 2025 57035 2275 58045 ;
    LAYER M1 ;
      RECT 2025 59135 2275 60145 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2455 35615 2705 39145 ;
    LAYER M1 ;
      RECT 2455 41495 2705 45025 ;
    LAYER M1 ;
      RECT 2455 47375 2705 50905 ;
    LAYER M1 ;
      RECT 2455 53255 2705 56785 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 15625 ;
    LAYER M1 ;
      RECT 2885 15875 3135 16885 ;
    LAYER M1 ;
      RECT 2885 17975 3135 21505 ;
    LAYER M1 ;
      RECT 2885 21755 3135 22765 ;
    LAYER M1 ;
      RECT 2885 23855 3135 27385 ;
    LAYER M1 ;
      RECT 2885 27635 3135 28645 ;
    LAYER M1 ;
      RECT 2885 29735 3135 33265 ;
    LAYER M1 ;
      RECT 2885 33515 3135 34525 ;
    LAYER M1 ;
      RECT 2885 35615 3135 39145 ;
    LAYER M1 ;
      RECT 2885 39395 3135 40405 ;
    LAYER M1 ;
      RECT 2885 41495 3135 45025 ;
    LAYER M1 ;
      RECT 2885 45275 3135 46285 ;
    LAYER M1 ;
      RECT 2885 47375 3135 50905 ;
    LAYER M1 ;
      RECT 2885 51155 3135 52165 ;
    LAYER M1 ;
      RECT 2885 53255 3135 56785 ;
    LAYER M1 ;
      RECT 2885 57035 3135 58045 ;
    LAYER M1 ;
      RECT 2885 59135 3135 60145 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 23855 3565 27385 ;
    LAYER M1 ;
      RECT 3315 29735 3565 33265 ;
    LAYER M1 ;
      RECT 3315 35615 3565 39145 ;
    LAYER M1 ;
      RECT 3315 41495 3565 45025 ;
    LAYER M1 ;
      RECT 3315 47375 3565 50905 ;
    LAYER M1 ;
      RECT 3315 53255 3565 56785 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 15625 ;
    LAYER M1 ;
      RECT 3745 15875 3995 16885 ;
    LAYER M1 ;
      RECT 3745 17975 3995 21505 ;
    LAYER M1 ;
      RECT 3745 21755 3995 22765 ;
    LAYER M1 ;
      RECT 3745 23855 3995 27385 ;
    LAYER M1 ;
      RECT 3745 27635 3995 28645 ;
    LAYER M1 ;
      RECT 3745 29735 3995 33265 ;
    LAYER M1 ;
      RECT 3745 33515 3995 34525 ;
    LAYER M1 ;
      RECT 3745 35615 3995 39145 ;
    LAYER M1 ;
      RECT 3745 39395 3995 40405 ;
    LAYER M1 ;
      RECT 3745 41495 3995 45025 ;
    LAYER M1 ;
      RECT 3745 45275 3995 46285 ;
    LAYER M1 ;
      RECT 3745 47375 3995 50905 ;
    LAYER M1 ;
      RECT 3745 51155 3995 52165 ;
    LAYER M1 ;
      RECT 3745 53255 3995 56785 ;
    LAYER M1 ;
      RECT 3745 57035 3995 58045 ;
    LAYER M1 ;
      RECT 3745 59135 3995 60145 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4175 17975 4425 21505 ;
    LAYER M1 ;
      RECT 4175 23855 4425 27385 ;
    LAYER M1 ;
      RECT 4175 29735 4425 33265 ;
    LAYER M1 ;
      RECT 4175 35615 4425 39145 ;
    LAYER M1 ;
      RECT 4175 41495 4425 45025 ;
    LAYER M1 ;
      RECT 4175 47375 4425 50905 ;
    LAYER M1 ;
      RECT 4175 53255 4425 56785 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 15625 ;
    LAYER M1 ;
      RECT 4605 15875 4855 16885 ;
    LAYER M1 ;
      RECT 4605 17975 4855 21505 ;
    LAYER M1 ;
      RECT 4605 21755 4855 22765 ;
    LAYER M1 ;
      RECT 4605 23855 4855 27385 ;
    LAYER M1 ;
      RECT 4605 27635 4855 28645 ;
    LAYER M1 ;
      RECT 4605 29735 4855 33265 ;
    LAYER M1 ;
      RECT 4605 33515 4855 34525 ;
    LAYER M1 ;
      RECT 4605 35615 4855 39145 ;
    LAYER M1 ;
      RECT 4605 39395 4855 40405 ;
    LAYER M1 ;
      RECT 4605 41495 4855 45025 ;
    LAYER M1 ;
      RECT 4605 45275 4855 46285 ;
    LAYER M1 ;
      RECT 4605 47375 4855 50905 ;
    LAYER M1 ;
      RECT 4605 51155 4855 52165 ;
    LAYER M1 ;
      RECT 4605 53255 4855 56785 ;
    LAYER M1 ;
      RECT 4605 57035 4855 58045 ;
    LAYER M1 ;
      RECT 4605 59135 4855 60145 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5035 12095 5285 15625 ;
    LAYER M1 ;
      RECT 5035 17975 5285 21505 ;
    LAYER M1 ;
      RECT 5035 23855 5285 27385 ;
    LAYER M1 ;
      RECT 5035 29735 5285 33265 ;
    LAYER M1 ;
      RECT 5035 35615 5285 39145 ;
    LAYER M1 ;
      RECT 5035 41495 5285 45025 ;
    LAYER M1 ;
      RECT 5035 47375 5285 50905 ;
    LAYER M1 ;
      RECT 5035 53255 5285 56785 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 15625 ;
    LAYER M1 ;
      RECT 5465 15875 5715 16885 ;
    LAYER M1 ;
      RECT 5465 17975 5715 21505 ;
    LAYER M1 ;
      RECT 5465 21755 5715 22765 ;
    LAYER M1 ;
      RECT 5465 23855 5715 27385 ;
    LAYER M1 ;
      RECT 5465 27635 5715 28645 ;
    LAYER M1 ;
      RECT 5465 29735 5715 33265 ;
    LAYER M1 ;
      RECT 5465 33515 5715 34525 ;
    LAYER M1 ;
      RECT 5465 35615 5715 39145 ;
    LAYER M1 ;
      RECT 5465 39395 5715 40405 ;
    LAYER M1 ;
      RECT 5465 41495 5715 45025 ;
    LAYER M1 ;
      RECT 5465 45275 5715 46285 ;
    LAYER M1 ;
      RECT 5465 47375 5715 50905 ;
    LAYER M1 ;
      RECT 5465 51155 5715 52165 ;
    LAYER M1 ;
      RECT 5465 53255 5715 56785 ;
    LAYER M1 ;
      RECT 5465 57035 5715 58045 ;
    LAYER M1 ;
      RECT 5465 59135 5715 60145 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 5895 12095 6145 15625 ;
    LAYER M1 ;
      RECT 5895 17975 6145 21505 ;
    LAYER M1 ;
      RECT 5895 23855 6145 27385 ;
    LAYER M1 ;
      RECT 5895 29735 6145 33265 ;
    LAYER M1 ;
      RECT 5895 35615 6145 39145 ;
    LAYER M1 ;
      RECT 5895 41495 6145 45025 ;
    LAYER M1 ;
      RECT 5895 47375 6145 50905 ;
    LAYER M1 ;
      RECT 5895 53255 6145 56785 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 9745 ;
    LAYER M1 ;
      RECT 6325 9995 6575 11005 ;
    LAYER M1 ;
      RECT 6325 12095 6575 15625 ;
    LAYER M1 ;
      RECT 6325 15875 6575 16885 ;
    LAYER M1 ;
      RECT 6325 17975 6575 21505 ;
    LAYER M1 ;
      RECT 6325 21755 6575 22765 ;
    LAYER M1 ;
      RECT 6325 23855 6575 27385 ;
    LAYER M1 ;
      RECT 6325 27635 6575 28645 ;
    LAYER M1 ;
      RECT 6325 29735 6575 33265 ;
    LAYER M1 ;
      RECT 6325 33515 6575 34525 ;
    LAYER M1 ;
      RECT 6325 35615 6575 39145 ;
    LAYER M1 ;
      RECT 6325 39395 6575 40405 ;
    LAYER M1 ;
      RECT 6325 41495 6575 45025 ;
    LAYER M1 ;
      RECT 6325 45275 6575 46285 ;
    LAYER M1 ;
      RECT 6325 47375 6575 50905 ;
    LAYER M1 ;
      RECT 6325 51155 6575 52165 ;
    LAYER M1 ;
      RECT 6325 53255 6575 56785 ;
    LAYER M1 ;
      RECT 6325 57035 6575 58045 ;
    LAYER M1 ;
      RECT 6325 59135 6575 60145 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 6215 7005 9745 ;
    LAYER M1 ;
      RECT 6755 12095 7005 15625 ;
    LAYER M1 ;
      RECT 6755 17975 7005 21505 ;
    LAYER M1 ;
      RECT 6755 23855 7005 27385 ;
    LAYER M1 ;
      RECT 6755 29735 7005 33265 ;
    LAYER M1 ;
      RECT 6755 35615 7005 39145 ;
    LAYER M1 ;
      RECT 6755 41495 7005 45025 ;
    LAYER M1 ;
      RECT 6755 47375 7005 50905 ;
    LAYER M1 ;
      RECT 6755 53255 7005 56785 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 9745 ;
    LAYER M1 ;
      RECT 7185 9995 7435 11005 ;
    LAYER M1 ;
      RECT 7185 12095 7435 15625 ;
    LAYER M1 ;
      RECT 7185 15875 7435 16885 ;
    LAYER M1 ;
      RECT 7185 17975 7435 21505 ;
    LAYER M1 ;
      RECT 7185 21755 7435 22765 ;
    LAYER M1 ;
      RECT 7185 23855 7435 27385 ;
    LAYER M1 ;
      RECT 7185 27635 7435 28645 ;
    LAYER M1 ;
      RECT 7185 29735 7435 33265 ;
    LAYER M1 ;
      RECT 7185 33515 7435 34525 ;
    LAYER M1 ;
      RECT 7185 35615 7435 39145 ;
    LAYER M1 ;
      RECT 7185 39395 7435 40405 ;
    LAYER M1 ;
      RECT 7185 41495 7435 45025 ;
    LAYER M1 ;
      RECT 7185 45275 7435 46285 ;
    LAYER M1 ;
      RECT 7185 47375 7435 50905 ;
    LAYER M1 ;
      RECT 7185 51155 7435 52165 ;
    LAYER M1 ;
      RECT 7185 53255 7435 56785 ;
    LAYER M1 ;
      RECT 7185 57035 7435 58045 ;
    LAYER M1 ;
      RECT 7185 59135 7435 60145 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 7615 6215 7865 9745 ;
    LAYER M1 ;
      RECT 7615 12095 7865 15625 ;
    LAYER M1 ;
      RECT 7615 17975 7865 21505 ;
    LAYER M1 ;
      RECT 7615 23855 7865 27385 ;
    LAYER M1 ;
      RECT 7615 29735 7865 33265 ;
    LAYER M1 ;
      RECT 7615 35615 7865 39145 ;
    LAYER M1 ;
      RECT 7615 41495 7865 45025 ;
    LAYER M1 ;
      RECT 7615 47375 7865 50905 ;
    LAYER M1 ;
      RECT 7615 53255 7865 56785 ;
    LAYER M2 ;
      RECT 1120 280 7480 560 ;
    LAYER M2 ;
      RECT 1120 4480 7480 4760 ;
    LAYER M2 ;
      RECT 690 700 7910 980 ;
    LAYER M2 ;
      RECT 1120 6160 7480 6440 ;
    LAYER M2 ;
      RECT 1120 10360 7480 10640 ;
    LAYER M2 ;
      RECT 690 6580 7910 6860 ;
    LAYER M2 ;
      RECT 1120 12040 7480 12320 ;
    LAYER M2 ;
      RECT 1120 16240 7480 16520 ;
    LAYER M2 ;
      RECT 690 12460 7910 12740 ;
    LAYER M2 ;
      RECT 1120 17920 7480 18200 ;
    LAYER M2 ;
      RECT 1120 22120 7480 22400 ;
    LAYER M2 ;
      RECT 690 18340 7910 18620 ;
    LAYER M2 ;
      RECT 1120 23800 7480 24080 ;
    LAYER M2 ;
      RECT 1120 28000 7480 28280 ;
    LAYER M2 ;
      RECT 690 24220 7910 24500 ;
    LAYER M2 ;
      RECT 1120 29680 7480 29960 ;
    LAYER M2 ;
      RECT 1120 33880 7480 34160 ;
    LAYER M2 ;
      RECT 690 30100 7910 30380 ;
    LAYER M2 ;
      RECT 1120 35560 7480 35840 ;
    LAYER M2 ;
      RECT 1120 39760 7480 40040 ;
    LAYER M2 ;
      RECT 690 35980 7910 36260 ;
    LAYER M2 ;
      RECT 1120 41440 7480 41720 ;
    LAYER M2 ;
      RECT 1120 45640 7480 45920 ;
    LAYER M2 ;
      RECT 690 41860 7910 42140 ;
    LAYER M2 ;
      RECT 1120 47320 7480 47600 ;
    LAYER M2 ;
      RECT 1120 51520 7480 51800 ;
    LAYER M2 ;
      RECT 690 47740 7910 48020 ;
    LAYER M2 ;
      RECT 1120 53200 7480 53480 ;
    LAYER M2 ;
      RECT 1120 57400 7480 57680 ;
    LAYER M2 ;
      RECT 1120 59500 7480 59780 ;
    LAYER M2 ;
      RECT 690 53620 7910 53900 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53255 1375 53425 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59555 1375 59725 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 29735 2235 29905 ;
    LAYER V1 ;
      RECT 2065 33935 2235 34105 ;
    LAYER V1 ;
      RECT 2065 35615 2235 35785 ;
    LAYER V1 ;
      RECT 2065 39815 2235 39985 ;
    LAYER V1 ;
      RECT 2065 41495 2235 41665 ;
    LAYER V1 ;
      RECT 2065 45695 2235 45865 ;
    LAYER V1 ;
      RECT 2065 47375 2235 47545 ;
    LAYER V1 ;
      RECT 2065 51575 2235 51745 ;
    LAYER V1 ;
      RECT 2065 53255 2235 53425 ;
    LAYER V1 ;
      RECT 2065 57455 2235 57625 ;
    LAYER V1 ;
      RECT 2065 59555 2235 59725 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12095 3095 12265 ;
    LAYER V1 ;
      RECT 2925 16295 3095 16465 ;
    LAYER V1 ;
      RECT 2925 17975 3095 18145 ;
    LAYER V1 ;
      RECT 2925 22175 3095 22345 ;
    LAYER V1 ;
      RECT 2925 23855 3095 24025 ;
    LAYER V1 ;
      RECT 2925 28055 3095 28225 ;
    LAYER V1 ;
      RECT 2925 29735 3095 29905 ;
    LAYER V1 ;
      RECT 2925 33935 3095 34105 ;
    LAYER V1 ;
      RECT 2925 35615 3095 35785 ;
    LAYER V1 ;
      RECT 2925 39815 3095 39985 ;
    LAYER V1 ;
      RECT 2925 41495 3095 41665 ;
    LAYER V1 ;
      RECT 2925 45695 3095 45865 ;
    LAYER V1 ;
      RECT 2925 47375 3095 47545 ;
    LAYER V1 ;
      RECT 2925 51575 3095 51745 ;
    LAYER V1 ;
      RECT 2925 53255 3095 53425 ;
    LAYER V1 ;
      RECT 2925 57455 3095 57625 ;
    LAYER V1 ;
      RECT 2925 59555 3095 59725 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12095 3955 12265 ;
    LAYER V1 ;
      RECT 3785 16295 3955 16465 ;
    LAYER V1 ;
      RECT 3785 17975 3955 18145 ;
    LAYER V1 ;
      RECT 3785 22175 3955 22345 ;
    LAYER V1 ;
      RECT 3785 23855 3955 24025 ;
    LAYER V1 ;
      RECT 3785 28055 3955 28225 ;
    LAYER V1 ;
      RECT 3785 29735 3955 29905 ;
    LAYER V1 ;
      RECT 3785 33935 3955 34105 ;
    LAYER V1 ;
      RECT 3785 35615 3955 35785 ;
    LAYER V1 ;
      RECT 3785 39815 3955 39985 ;
    LAYER V1 ;
      RECT 3785 41495 3955 41665 ;
    LAYER V1 ;
      RECT 3785 45695 3955 45865 ;
    LAYER V1 ;
      RECT 3785 47375 3955 47545 ;
    LAYER V1 ;
      RECT 3785 51575 3955 51745 ;
    LAYER V1 ;
      RECT 3785 53255 3955 53425 ;
    LAYER V1 ;
      RECT 3785 57455 3955 57625 ;
    LAYER V1 ;
      RECT 3785 59555 3955 59725 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12095 4815 12265 ;
    LAYER V1 ;
      RECT 4645 16295 4815 16465 ;
    LAYER V1 ;
      RECT 4645 17975 4815 18145 ;
    LAYER V1 ;
      RECT 4645 22175 4815 22345 ;
    LAYER V1 ;
      RECT 4645 23855 4815 24025 ;
    LAYER V1 ;
      RECT 4645 28055 4815 28225 ;
    LAYER V1 ;
      RECT 4645 29735 4815 29905 ;
    LAYER V1 ;
      RECT 4645 33935 4815 34105 ;
    LAYER V1 ;
      RECT 4645 35615 4815 35785 ;
    LAYER V1 ;
      RECT 4645 39815 4815 39985 ;
    LAYER V1 ;
      RECT 4645 41495 4815 41665 ;
    LAYER V1 ;
      RECT 4645 45695 4815 45865 ;
    LAYER V1 ;
      RECT 4645 47375 4815 47545 ;
    LAYER V1 ;
      RECT 4645 51575 4815 51745 ;
    LAYER V1 ;
      RECT 4645 53255 4815 53425 ;
    LAYER V1 ;
      RECT 4645 57455 4815 57625 ;
    LAYER V1 ;
      RECT 4645 59555 4815 59725 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12095 5675 12265 ;
    LAYER V1 ;
      RECT 5505 16295 5675 16465 ;
    LAYER V1 ;
      RECT 5505 17975 5675 18145 ;
    LAYER V1 ;
      RECT 5505 22175 5675 22345 ;
    LAYER V1 ;
      RECT 5505 23855 5675 24025 ;
    LAYER V1 ;
      RECT 5505 28055 5675 28225 ;
    LAYER V1 ;
      RECT 5505 29735 5675 29905 ;
    LAYER V1 ;
      RECT 5505 33935 5675 34105 ;
    LAYER V1 ;
      RECT 5505 35615 5675 35785 ;
    LAYER V1 ;
      RECT 5505 39815 5675 39985 ;
    LAYER V1 ;
      RECT 5505 41495 5675 41665 ;
    LAYER V1 ;
      RECT 5505 45695 5675 45865 ;
    LAYER V1 ;
      RECT 5505 47375 5675 47545 ;
    LAYER V1 ;
      RECT 5505 51575 5675 51745 ;
    LAYER V1 ;
      RECT 5505 53255 5675 53425 ;
    LAYER V1 ;
      RECT 5505 57455 5675 57625 ;
    LAYER V1 ;
      RECT 5505 59555 5675 59725 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6215 6535 6385 ;
    LAYER V1 ;
      RECT 6365 10415 6535 10585 ;
    LAYER V1 ;
      RECT 6365 12095 6535 12265 ;
    LAYER V1 ;
      RECT 6365 16295 6535 16465 ;
    LAYER V1 ;
      RECT 6365 17975 6535 18145 ;
    LAYER V1 ;
      RECT 6365 22175 6535 22345 ;
    LAYER V1 ;
      RECT 6365 23855 6535 24025 ;
    LAYER V1 ;
      RECT 6365 28055 6535 28225 ;
    LAYER V1 ;
      RECT 6365 29735 6535 29905 ;
    LAYER V1 ;
      RECT 6365 33935 6535 34105 ;
    LAYER V1 ;
      RECT 6365 35615 6535 35785 ;
    LAYER V1 ;
      RECT 6365 39815 6535 39985 ;
    LAYER V1 ;
      RECT 6365 41495 6535 41665 ;
    LAYER V1 ;
      RECT 6365 45695 6535 45865 ;
    LAYER V1 ;
      RECT 6365 47375 6535 47545 ;
    LAYER V1 ;
      RECT 6365 51575 6535 51745 ;
    LAYER V1 ;
      RECT 6365 53255 6535 53425 ;
    LAYER V1 ;
      RECT 6365 57455 6535 57625 ;
    LAYER V1 ;
      RECT 6365 59555 6535 59725 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6215 7395 6385 ;
    LAYER V1 ;
      RECT 7225 10415 7395 10585 ;
    LAYER V1 ;
      RECT 7225 12095 7395 12265 ;
    LAYER V1 ;
      RECT 7225 16295 7395 16465 ;
    LAYER V1 ;
      RECT 7225 17975 7395 18145 ;
    LAYER V1 ;
      RECT 7225 22175 7395 22345 ;
    LAYER V1 ;
      RECT 7225 23855 7395 24025 ;
    LAYER V1 ;
      RECT 7225 28055 7395 28225 ;
    LAYER V1 ;
      RECT 7225 29735 7395 29905 ;
    LAYER V1 ;
      RECT 7225 33935 7395 34105 ;
    LAYER V1 ;
      RECT 7225 35615 7395 35785 ;
    LAYER V1 ;
      RECT 7225 39815 7395 39985 ;
    LAYER V1 ;
      RECT 7225 41495 7395 41665 ;
    LAYER V1 ;
      RECT 7225 45695 7395 45865 ;
    LAYER V1 ;
      RECT 7225 47375 7395 47545 ;
    LAYER V1 ;
      RECT 7225 51575 7395 51745 ;
    LAYER V1 ;
      RECT 7225 53255 7395 53425 ;
    LAYER V1 ;
      RECT 7225 57455 7395 57625 ;
    LAYER V1 ;
      RECT 7225 59555 7395 59725 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 775 53675 945 53845 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 1635 53675 1805 53845 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 2495 30155 2665 30325 ;
    LAYER V1 ;
      RECT 2495 36035 2665 36205 ;
    LAYER V1 ;
      RECT 2495 41915 2665 42085 ;
    LAYER V1 ;
      RECT 2495 47795 2665 47965 ;
    LAYER V1 ;
      RECT 2495 53675 2665 53845 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 18395 3525 18565 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 3355 30155 3525 30325 ;
    LAYER V1 ;
      RECT 3355 36035 3525 36205 ;
    LAYER V1 ;
      RECT 3355 41915 3525 42085 ;
    LAYER V1 ;
      RECT 3355 47795 3525 47965 ;
    LAYER V1 ;
      RECT 3355 53675 3525 53845 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 4215 12515 4385 12685 ;
    LAYER V1 ;
      RECT 4215 18395 4385 18565 ;
    LAYER V1 ;
      RECT 4215 24275 4385 24445 ;
    LAYER V1 ;
      RECT 4215 30155 4385 30325 ;
    LAYER V1 ;
      RECT 4215 36035 4385 36205 ;
    LAYER V1 ;
      RECT 4215 41915 4385 42085 ;
    LAYER V1 ;
      RECT 4215 47795 4385 47965 ;
    LAYER V1 ;
      RECT 4215 53675 4385 53845 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 5075 12515 5245 12685 ;
    LAYER V1 ;
      RECT 5075 18395 5245 18565 ;
    LAYER V1 ;
      RECT 5075 24275 5245 24445 ;
    LAYER V1 ;
      RECT 5075 30155 5245 30325 ;
    LAYER V1 ;
      RECT 5075 36035 5245 36205 ;
    LAYER V1 ;
      RECT 5075 41915 5245 42085 ;
    LAYER V1 ;
      RECT 5075 47795 5245 47965 ;
    LAYER V1 ;
      RECT 5075 53675 5245 53845 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 5935 6635 6105 6805 ;
    LAYER V1 ;
      RECT 5935 12515 6105 12685 ;
    LAYER V1 ;
      RECT 5935 18395 6105 18565 ;
    LAYER V1 ;
      RECT 5935 24275 6105 24445 ;
    LAYER V1 ;
      RECT 5935 30155 6105 30325 ;
    LAYER V1 ;
      RECT 5935 36035 6105 36205 ;
    LAYER V1 ;
      RECT 5935 41915 6105 42085 ;
    LAYER V1 ;
      RECT 5935 47795 6105 47965 ;
    LAYER V1 ;
      RECT 5935 53675 6105 53845 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 6795 12515 6965 12685 ;
    LAYER V1 ;
      RECT 6795 18395 6965 18565 ;
    LAYER V1 ;
      RECT 6795 24275 6965 24445 ;
    LAYER V1 ;
      RECT 6795 30155 6965 30325 ;
    LAYER V1 ;
      RECT 6795 36035 6965 36205 ;
    LAYER V1 ;
      RECT 6795 41915 6965 42085 ;
    LAYER V1 ;
      RECT 6795 47795 6965 47965 ;
    LAYER V1 ;
      RECT 6795 53675 6965 53845 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 7655 6635 7825 6805 ;
    LAYER V1 ;
      RECT 7655 12515 7825 12685 ;
    LAYER V1 ;
      RECT 7655 18395 7825 18565 ;
    LAYER V1 ;
      RECT 7655 24275 7825 24445 ;
    LAYER V1 ;
      RECT 7655 30155 7825 30325 ;
    LAYER V1 ;
      RECT 7655 36035 7825 36205 ;
    LAYER V1 ;
      RECT 7655 41915 7825 42085 ;
    LAYER V1 ;
      RECT 7655 47795 7825 47965 ;
    LAYER V1 ;
      RECT 7655 53675 7825 53845 ;
    LAYER V2 ;
      RECT 3795 345 3945 495 ;
    LAYER V2 ;
      RECT 3795 6225 3945 6375 ;
    LAYER V2 ;
      RECT 3795 12105 3945 12255 ;
    LAYER V2 ;
      RECT 3795 17985 3945 18135 ;
    LAYER V2 ;
      RECT 3795 23865 3945 24015 ;
    LAYER V2 ;
      RECT 3795 29745 3945 29895 ;
    LAYER V2 ;
      RECT 3795 35625 3945 35775 ;
    LAYER V2 ;
      RECT 3795 41505 3945 41655 ;
    LAYER V2 ;
      RECT 3795 47385 3945 47535 ;
    LAYER V2 ;
      RECT 3795 53265 3945 53415 ;
    LAYER V2 ;
      RECT 4225 4545 4375 4695 ;
    LAYER V2 ;
      RECT 4225 10425 4375 10575 ;
    LAYER V2 ;
      RECT 4225 16305 4375 16455 ;
    LAYER V2 ;
      RECT 4225 22185 4375 22335 ;
    LAYER V2 ;
      RECT 4225 28065 4375 28215 ;
    LAYER V2 ;
      RECT 4225 33945 4375 34095 ;
    LAYER V2 ;
      RECT 4225 39825 4375 39975 ;
    LAYER V2 ;
      RECT 4225 45705 4375 45855 ;
    LAYER V2 ;
      RECT 4225 51585 4375 51735 ;
    LAYER V2 ;
      RECT 4225 57465 4375 57615 ;
    LAYER V2 ;
      RECT 4655 765 4805 915 ;
    LAYER V2 ;
      RECT 4655 6645 4805 6795 ;
    LAYER V2 ;
      RECT 4655 12525 4805 12675 ;
    LAYER V2 ;
      RECT 4655 18405 4805 18555 ;
    LAYER V2 ;
      RECT 4655 24285 4805 24435 ;
    LAYER V2 ;
      RECT 4655 30165 4805 30315 ;
    LAYER V2 ;
      RECT 4655 36045 4805 36195 ;
    LAYER V2 ;
      RECT 4655 41925 4805 42075 ;
    LAYER V2 ;
      RECT 4655 47805 4805 47955 ;
    LAYER V2 ;
      RECT 4655 53685 4805 53835 ;
    LAYER V2 ;
      RECT 4655 59565 4805 59715 ;
  END
END NMOS_S_80601593_X8_Y10
