MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 67.67 BY 56.87 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 28.24 0.26 28.52 28.3 ;
      LAYER M3 ;
        RECT 38.56 4.46 38.84 28.3 ;
      LAYER M3 ;
        RECT 28.24 14.935 28.52 15.305 ;
      LAYER M2 ;
        RECT 28.38 14.98 38.7 15.26 ;
      LAYER M3 ;
        RECT 38.56 14.935 38.84 15.305 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 51.89 24.62 52.17 30.82 ;
      LAYER M3 ;
        RECT 50.6 31.34 50.88 49.3 ;
      LAYER M3 ;
        RECT 51.89 30.66 52.17 31.5 ;
      LAYER M4 ;
        RECT 50.74 31.1 52.03 31.9 ;
      LAYER M3 ;
        RECT 50.6 31.315 50.88 31.685 ;
    END
  END VOUT
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 11.2 22.1 11.48 ;
    END
  END VINN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 44.98 11.2 65.96 11.48 ;
    END
  END VINP
  OBS 
  LAYER M3 ;
        RECT 14.91 24.62 15.19 30.82 ;
  LAYER M3 ;
        RECT 16.63 31.34 16.91 53.5 ;
  LAYER M3 ;
        RECT 50.17 35.54 50.45 53.5 ;
  LAYER M3 ;
        RECT 14.91 30.66 15.19 31.5 ;
  LAYER M4 ;
        RECT 15.05 31.1 16.77 31.9 ;
  LAYER M3 ;
        RECT 16.63 31.315 16.91 31.685 ;
  LAYER M3 ;
        RECT 16.63 37.615 16.91 37.985 ;
  LAYER M4 ;
        RECT 16.77 37.4 50.31 38.2 ;
  LAYER M3 ;
        RECT 50.17 37.615 50.45 37.985 ;
  LAYER M3 ;
        RECT 14.91 31.315 15.19 31.685 ;
  LAYER M4 ;
        RECT 14.885 31.1 15.215 31.9 ;
  LAYER M3 ;
        RECT 16.63 31.315 16.91 31.685 ;
  LAYER M4 ;
        RECT 16.605 31.1 16.935 31.9 ;
  LAYER M3 ;
        RECT 14.91 31.315 15.19 31.685 ;
  LAYER M4 ;
        RECT 14.885 31.1 15.215 31.9 ;
  LAYER M3 ;
        RECT 16.63 31.315 16.91 31.685 ;
  LAYER M4 ;
        RECT 16.605 31.1 16.935 31.9 ;
  LAYER M3 ;
        RECT 14.91 31.315 15.19 31.685 ;
  LAYER M4 ;
        RECT 14.885 31.1 15.215 31.9 ;
  LAYER M3 ;
        RECT 16.63 31.315 16.91 31.685 ;
  LAYER M4 ;
        RECT 16.605 31.1 16.935 31.9 ;
  LAYER M3 ;
        RECT 16.63 37.615 16.91 37.985 ;
  LAYER M4 ;
        RECT 16.605 37.4 16.935 38.2 ;
  LAYER M3 ;
        RECT 50.17 37.615 50.45 37.985 ;
  LAYER M4 ;
        RECT 50.145 37.4 50.475 38.2 ;
  LAYER M3 ;
        RECT 14.91 31.315 15.19 31.685 ;
  LAYER M4 ;
        RECT 14.885 31.1 15.215 31.9 ;
  LAYER M3 ;
        RECT 16.63 31.315 16.91 31.685 ;
  LAYER M4 ;
        RECT 16.605 31.1 16.935 31.9 ;
  LAYER M3 ;
        RECT 16.63 37.615 16.91 37.985 ;
  LAYER M4 ;
        RECT 16.605 37.4 16.935 38.2 ;
  LAYER M3 ;
        RECT 50.17 37.615 50.45 37.985 ;
  LAYER M4 ;
        RECT 50.145 37.4 50.475 38.2 ;
  LAYER M3 ;
        RECT 2.01 16.22 2.29 26.62 ;
  LAYER M3 ;
        RECT 14.48 20.42 14.76 26.62 ;
  LAYER M2 ;
        RECT 1.12 15.4 22.1 15.68 ;
  LAYER M3 ;
        RECT 2.01 20.815 2.29 21.185 ;
  LAYER M2 ;
        RECT 2.15 20.86 14.62 21.14 ;
  LAYER M3 ;
        RECT 14.48 20.815 14.76 21.185 ;
  LAYER M3 ;
        RECT 2.01 15.54 2.29 16.38 ;
  LAYER M2 ;
        RECT 1.99 15.4 2.31 15.68 ;
  LAYER M2 ;
        RECT 1.99 20.86 2.31 21.14 ;
  LAYER M3 ;
        RECT 2.01 20.84 2.29 21.16 ;
  LAYER M2 ;
        RECT 14.46 20.86 14.78 21.14 ;
  LAYER M3 ;
        RECT 14.48 20.84 14.76 21.16 ;
  LAYER M2 ;
        RECT 1.99 20.86 2.31 21.14 ;
  LAYER M3 ;
        RECT 2.01 20.84 2.29 21.16 ;
  LAYER M2 ;
        RECT 14.46 20.86 14.78 21.14 ;
  LAYER M3 ;
        RECT 14.48 20.84 14.76 21.16 ;
  LAYER M2 ;
        RECT 1.99 15.4 2.31 15.68 ;
  LAYER M3 ;
        RECT 2.01 15.38 2.29 15.7 ;
  LAYER M2 ;
        RECT 1.99 20.86 2.31 21.14 ;
  LAYER M3 ;
        RECT 2.01 20.84 2.29 21.16 ;
  LAYER M2 ;
        RECT 14.46 20.86 14.78 21.14 ;
  LAYER M3 ;
        RECT 14.48 20.84 14.76 21.16 ;
  LAYER M2 ;
        RECT 1.99 15.4 2.31 15.68 ;
  LAYER M3 ;
        RECT 2.01 15.38 2.29 15.7 ;
  LAYER M2 ;
        RECT 1.99 20.86 2.31 21.14 ;
  LAYER M3 ;
        RECT 2.01 20.84 2.29 21.16 ;
  LAYER M2 ;
        RECT 14.46 20.86 14.78 21.14 ;
  LAYER M3 ;
        RECT 14.48 20.84 14.76 21.16 ;
  LAYER M2 ;
        RECT 44.98 15.4 65.96 15.68 ;
  LAYER M3 ;
        RECT 52.32 20.42 52.6 26.62 ;
  LAYER M3 ;
        RECT 64.79 16.22 65.07 26.62 ;
  LAYER M2 ;
        RECT 52.3 15.4 52.62 15.68 ;
  LAYER M3 ;
        RECT 52.32 15.54 52.6 20.58 ;
  LAYER M2 ;
        RECT 64.77 15.4 65.09 15.68 ;
  LAYER M3 ;
        RECT 64.79 15.54 65.07 16.38 ;
  LAYER M2 ;
        RECT 52.3 15.4 52.62 15.68 ;
  LAYER M3 ;
        RECT 52.32 15.38 52.6 15.7 ;
  LAYER M2 ;
        RECT 52.3 15.4 52.62 15.68 ;
  LAYER M3 ;
        RECT 52.32 15.38 52.6 15.7 ;
  LAYER M2 ;
        RECT 52.3 15.4 52.62 15.68 ;
  LAYER M3 ;
        RECT 52.32 15.38 52.6 15.7 ;
  LAYER M2 ;
        RECT 64.77 15.4 65.09 15.68 ;
  LAYER M3 ;
        RECT 64.79 15.38 65.07 15.7 ;
  LAYER M2 ;
        RECT 52.3 15.4 52.62 15.68 ;
  LAYER M3 ;
        RECT 52.32 15.38 52.6 15.7 ;
  LAYER M2 ;
        RECT 64.77 15.4 65.09 15.68 ;
  LAYER M3 ;
        RECT 64.79 15.38 65.07 15.7 ;
  LAYER M2 ;
        RECT 0.69 14.98 22.53 15.26 ;
  LAYER M3 ;
        RECT 38.13 0.26 38.41 24.1 ;
  LAYER M2 ;
        RECT 44.55 14.98 66.39 15.26 ;
  LAYER M2 ;
        RECT 22.36 14.98 25.8 15.26 ;
  LAYER M3 ;
        RECT 25.66 14.7 25.94 15.12 ;
  LAYER M2 ;
        RECT 25.8 14.56 38.27 14.84 ;
  LAYER M3 ;
        RECT 38.13 14.515 38.41 14.885 ;
  LAYER M3 ;
        RECT 38.13 14.935 38.41 15.305 ;
  LAYER M4 ;
        RECT 38.27 14.72 39.56 15.52 ;
  LAYER M3 ;
        RECT 39.42 14.999 39.7 15.241 ;
  LAYER M2 ;
        RECT 39.56 14.98 44.72 15.26 ;
  LAYER M2 ;
        RECT 25.64 14.56 25.96 14.84 ;
  LAYER M3 ;
        RECT 25.66 14.54 25.94 14.86 ;
  LAYER M2 ;
        RECT 25.64 14.98 25.96 15.26 ;
  LAYER M3 ;
        RECT 25.66 14.96 25.94 15.28 ;
  LAYER M2 ;
        RECT 38.11 14.56 38.43 14.84 ;
  LAYER M3 ;
        RECT 38.13 14.54 38.41 14.86 ;
  LAYER M2 ;
        RECT 25.64 14.56 25.96 14.84 ;
  LAYER M3 ;
        RECT 25.66 14.54 25.94 14.86 ;
  LAYER M2 ;
        RECT 25.64 14.98 25.96 15.26 ;
  LAYER M3 ;
        RECT 25.66 14.96 25.94 15.28 ;
  LAYER M2 ;
        RECT 38.11 14.56 38.43 14.84 ;
  LAYER M3 ;
        RECT 38.13 14.54 38.41 14.86 ;
  LAYER M2 ;
        RECT 25.64 14.56 25.96 14.84 ;
  LAYER M3 ;
        RECT 25.66 14.54 25.94 14.86 ;
  LAYER M2 ;
        RECT 25.64 14.98 25.96 15.26 ;
  LAYER M3 ;
        RECT 25.66 14.96 25.94 15.28 ;
  LAYER M2 ;
        RECT 38.11 14.56 38.43 14.84 ;
  LAYER M3 ;
        RECT 38.13 14.54 38.41 14.86 ;
  LAYER M2 ;
        RECT 39.4 14.98 39.72 15.26 ;
  LAYER M3 ;
        RECT 39.42 14.96 39.7 15.28 ;
  LAYER M3 ;
        RECT 38.13 14.935 38.41 15.305 ;
  LAYER M4 ;
        RECT 38.105 14.72 38.435 15.52 ;
  LAYER M3 ;
        RECT 39.42 14.935 39.7 15.305 ;
  LAYER M4 ;
        RECT 39.395 14.72 39.725 15.52 ;
  LAYER M2 ;
        RECT 25.64 14.56 25.96 14.84 ;
  LAYER M3 ;
        RECT 25.66 14.54 25.94 14.86 ;
  LAYER M2 ;
        RECT 25.64 14.98 25.96 15.26 ;
  LAYER M3 ;
        RECT 25.66 14.96 25.94 15.28 ;
  LAYER M2 ;
        RECT 38.11 14.56 38.43 14.84 ;
  LAYER M3 ;
        RECT 38.13 14.54 38.41 14.86 ;
  LAYER M3 ;
        RECT 38.13 14.935 38.41 15.305 ;
  LAYER M4 ;
        RECT 38.105 14.72 38.435 15.52 ;
  LAYER M1 ;
        RECT 32.125 0.335 32.375 3.865 ;
  LAYER M1 ;
        RECT 32.125 4.115 32.375 5.125 ;
  LAYER M1 ;
        RECT 32.125 6.215 32.375 9.745 ;
  LAYER M1 ;
        RECT 32.125 9.995 32.375 11.005 ;
  LAYER M1 ;
        RECT 32.125 12.095 32.375 15.625 ;
  LAYER M1 ;
        RECT 32.125 15.875 32.375 16.885 ;
  LAYER M1 ;
        RECT 32.125 17.975 32.375 21.505 ;
  LAYER M1 ;
        RECT 32.125 21.755 32.375 22.765 ;
  LAYER M1 ;
        RECT 32.125 23.855 32.375 27.385 ;
  LAYER M1 ;
        RECT 32.125 27.635 32.375 28.645 ;
  LAYER M1 ;
        RECT 32.125 29.735 32.375 30.745 ;
  LAYER M1 ;
        RECT 32.555 0.335 32.805 3.865 ;
  LAYER M1 ;
        RECT 32.555 6.215 32.805 9.745 ;
  LAYER M1 ;
        RECT 32.555 12.095 32.805 15.625 ;
  LAYER M1 ;
        RECT 32.555 17.975 32.805 21.505 ;
  LAYER M1 ;
        RECT 32.555 23.855 32.805 27.385 ;
  LAYER M1 ;
        RECT 31.695 0.335 31.945 3.865 ;
  LAYER M1 ;
        RECT 31.695 6.215 31.945 9.745 ;
  LAYER M1 ;
        RECT 31.695 12.095 31.945 15.625 ;
  LAYER M1 ;
        RECT 31.695 17.975 31.945 21.505 ;
  LAYER M1 ;
        RECT 31.695 23.855 31.945 27.385 ;
  LAYER M1 ;
        RECT 31.265 0.335 31.515 3.865 ;
  LAYER M1 ;
        RECT 31.265 4.115 31.515 5.125 ;
  LAYER M1 ;
        RECT 31.265 6.215 31.515 9.745 ;
  LAYER M1 ;
        RECT 31.265 9.995 31.515 11.005 ;
  LAYER M1 ;
        RECT 31.265 12.095 31.515 15.625 ;
  LAYER M1 ;
        RECT 31.265 15.875 31.515 16.885 ;
  LAYER M1 ;
        RECT 31.265 17.975 31.515 21.505 ;
  LAYER M1 ;
        RECT 31.265 21.755 31.515 22.765 ;
  LAYER M1 ;
        RECT 31.265 23.855 31.515 27.385 ;
  LAYER M1 ;
        RECT 31.265 27.635 31.515 28.645 ;
  LAYER M1 ;
        RECT 31.265 29.735 31.515 30.745 ;
  LAYER M1 ;
        RECT 30.835 0.335 31.085 3.865 ;
  LAYER M1 ;
        RECT 30.835 6.215 31.085 9.745 ;
  LAYER M1 ;
        RECT 30.835 12.095 31.085 15.625 ;
  LAYER M1 ;
        RECT 30.835 17.975 31.085 21.505 ;
  LAYER M1 ;
        RECT 30.835 23.855 31.085 27.385 ;
  LAYER M1 ;
        RECT 30.405 0.335 30.655 3.865 ;
  LAYER M1 ;
        RECT 30.405 4.115 30.655 5.125 ;
  LAYER M1 ;
        RECT 30.405 6.215 30.655 9.745 ;
  LAYER M1 ;
        RECT 30.405 9.995 30.655 11.005 ;
  LAYER M1 ;
        RECT 30.405 12.095 30.655 15.625 ;
  LAYER M1 ;
        RECT 30.405 15.875 30.655 16.885 ;
  LAYER M1 ;
        RECT 30.405 17.975 30.655 21.505 ;
  LAYER M1 ;
        RECT 30.405 21.755 30.655 22.765 ;
  LAYER M1 ;
        RECT 30.405 23.855 30.655 27.385 ;
  LAYER M1 ;
        RECT 30.405 27.635 30.655 28.645 ;
  LAYER M1 ;
        RECT 30.405 29.735 30.655 30.745 ;
  LAYER M1 ;
        RECT 29.975 0.335 30.225 3.865 ;
  LAYER M1 ;
        RECT 29.975 6.215 30.225 9.745 ;
  LAYER M1 ;
        RECT 29.975 12.095 30.225 15.625 ;
  LAYER M1 ;
        RECT 29.975 17.975 30.225 21.505 ;
  LAYER M1 ;
        RECT 29.975 23.855 30.225 27.385 ;
  LAYER M1 ;
        RECT 29.545 0.335 29.795 3.865 ;
  LAYER M1 ;
        RECT 29.545 4.115 29.795 5.125 ;
  LAYER M1 ;
        RECT 29.545 6.215 29.795 9.745 ;
  LAYER M1 ;
        RECT 29.545 9.995 29.795 11.005 ;
  LAYER M1 ;
        RECT 29.545 12.095 29.795 15.625 ;
  LAYER M1 ;
        RECT 29.545 15.875 29.795 16.885 ;
  LAYER M1 ;
        RECT 29.545 17.975 29.795 21.505 ;
  LAYER M1 ;
        RECT 29.545 21.755 29.795 22.765 ;
  LAYER M1 ;
        RECT 29.545 23.855 29.795 27.385 ;
  LAYER M1 ;
        RECT 29.545 27.635 29.795 28.645 ;
  LAYER M1 ;
        RECT 29.545 29.735 29.795 30.745 ;
  LAYER M1 ;
        RECT 29.115 0.335 29.365 3.865 ;
  LAYER M1 ;
        RECT 29.115 6.215 29.365 9.745 ;
  LAYER M1 ;
        RECT 29.115 12.095 29.365 15.625 ;
  LAYER M1 ;
        RECT 29.115 17.975 29.365 21.505 ;
  LAYER M1 ;
        RECT 29.115 23.855 29.365 27.385 ;
  LAYER M1 ;
        RECT 28.685 0.335 28.935 3.865 ;
  LAYER M1 ;
        RECT 28.685 4.115 28.935 5.125 ;
  LAYER M1 ;
        RECT 28.685 6.215 28.935 9.745 ;
  LAYER M1 ;
        RECT 28.685 9.995 28.935 11.005 ;
  LAYER M1 ;
        RECT 28.685 12.095 28.935 15.625 ;
  LAYER M1 ;
        RECT 28.685 15.875 28.935 16.885 ;
  LAYER M1 ;
        RECT 28.685 17.975 28.935 21.505 ;
  LAYER M1 ;
        RECT 28.685 21.755 28.935 22.765 ;
  LAYER M1 ;
        RECT 28.685 23.855 28.935 27.385 ;
  LAYER M1 ;
        RECT 28.685 27.635 28.935 28.645 ;
  LAYER M1 ;
        RECT 28.685 29.735 28.935 30.745 ;
  LAYER M1 ;
        RECT 28.255 0.335 28.505 3.865 ;
  LAYER M1 ;
        RECT 28.255 6.215 28.505 9.745 ;
  LAYER M1 ;
        RECT 28.255 12.095 28.505 15.625 ;
  LAYER M1 ;
        RECT 28.255 17.975 28.505 21.505 ;
  LAYER M1 ;
        RECT 28.255 23.855 28.505 27.385 ;
  LAYER M1 ;
        RECT 27.825 0.335 28.075 3.865 ;
  LAYER M1 ;
        RECT 27.825 4.115 28.075 5.125 ;
  LAYER M1 ;
        RECT 27.825 6.215 28.075 9.745 ;
  LAYER M1 ;
        RECT 27.825 9.995 28.075 11.005 ;
  LAYER M1 ;
        RECT 27.825 12.095 28.075 15.625 ;
  LAYER M1 ;
        RECT 27.825 15.875 28.075 16.885 ;
  LAYER M1 ;
        RECT 27.825 17.975 28.075 21.505 ;
  LAYER M1 ;
        RECT 27.825 21.755 28.075 22.765 ;
  LAYER M1 ;
        RECT 27.825 23.855 28.075 27.385 ;
  LAYER M1 ;
        RECT 27.825 27.635 28.075 28.645 ;
  LAYER M1 ;
        RECT 27.825 29.735 28.075 30.745 ;
  LAYER M1 ;
        RECT 27.395 0.335 27.645 3.865 ;
  LAYER M1 ;
        RECT 27.395 6.215 27.645 9.745 ;
  LAYER M1 ;
        RECT 27.395 12.095 27.645 15.625 ;
  LAYER M1 ;
        RECT 27.395 17.975 27.645 21.505 ;
  LAYER M1 ;
        RECT 27.395 23.855 27.645 27.385 ;
  LAYER M1 ;
        RECT 26.965 0.335 27.215 3.865 ;
  LAYER M1 ;
        RECT 26.965 4.115 27.215 5.125 ;
  LAYER M1 ;
        RECT 26.965 6.215 27.215 9.745 ;
  LAYER M1 ;
        RECT 26.965 9.995 27.215 11.005 ;
  LAYER M1 ;
        RECT 26.965 12.095 27.215 15.625 ;
  LAYER M1 ;
        RECT 26.965 15.875 27.215 16.885 ;
  LAYER M1 ;
        RECT 26.965 17.975 27.215 21.505 ;
  LAYER M1 ;
        RECT 26.965 21.755 27.215 22.765 ;
  LAYER M1 ;
        RECT 26.965 23.855 27.215 27.385 ;
  LAYER M1 ;
        RECT 26.965 27.635 27.215 28.645 ;
  LAYER M1 ;
        RECT 26.965 29.735 27.215 30.745 ;
  LAYER M1 ;
        RECT 26.535 0.335 26.785 3.865 ;
  LAYER M1 ;
        RECT 26.535 6.215 26.785 9.745 ;
  LAYER M1 ;
        RECT 26.535 12.095 26.785 15.625 ;
  LAYER M1 ;
        RECT 26.535 17.975 26.785 21.505 ;
  LAYER M1 ;
        RECT 26.535 23.855 26.785 27.385 ;
  LAYER M1 ;
        RECT 26.105 0.335 26.355 3.865 ;
  LAYER M1 ;
        RECT 26.105 4.115 26.355 5.125 ;
  LAYER M1 ;
        RECT 26.105 6.215 26.355 9.745 ;
  LAYER M1 ;
        RECT 26.105 9.995 26.355 11.005 ;
  LAYER M1 ;
        RECT 26.105 12.095 26.355 15.625 ;
  LAYER M1 ;
        RECT 26.105 15.875 26.355 16.885 ;
  LAYER M1 ;
        RECT 26.105 17.975 26.355 21.505 ;
  LAYER M1 ;
        RECT 26.105 21.755 26.355 22.765 ;
  LAYER M1 ;
        RECT 26.105 23.855 26.355 27.385 ;
  LAYER M1 ;
        RECT 26.105 27.635 26.355 28.645 ;
  LAYER M1 ;
        RECT 26.105 29.735 26.355 30.745 ;
  LAYER M1 ;
        RECT 25.675 0.335 25.925 3.865 ;
  LAYER M1 ;
        RECT 25.675 6.215 25.925 9.745 ;
  LAYER M1 ;
        RECT 25.675 12.095 25.925 15.625 ;
  LAYER M1 ;
        RECT 25.675 17.975 25.925 21.505 ;
  LAYER M1 ;
        RECT 25.675 23.855 25.925 27.385 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 3.865 ;
  LAYER M1 ;
        RECT 25.245 4.115 25.495 5.125 ;
  LAYER M1 ;
        RECT 25.245 6.215 25.495 9.745 ;
  LAYER M1 ;
        RECT 25.245 9.995 25.495 11.005 ;
  LAYER M1 ;
        RECT 25.245 12.095 25.495 15.625 ;
  LAYER M1 ;
        RECT 25.245 15.875 25.495 16.885 ;
  LAYER M1 ;
        RECT 25.245 17.975 25.495 21.505 ;
  LAYER M1 ;
        RECT 25.245 21.755 25.495 22.765 ;
  LAYER M1 ;
        RECT 25.245 23.855 25.495 27.385 ;
  LAYER M1 ;
        RECT 25.245 27.635 25.495 28.645 ;
  LAYER M1 ;
        RECT 25.245 29.735 25.495 30.745 ;
  LAYER M1 ;
        RECT 24.815 0.335 25.065 3.865 ;
  LAYER M1 ;
        RECT 24.815 6.215 25.065 9.745 ;
  LAYER M1 ;
        RECT 24.815 12.095 25.065 15.625 ;
  LAYER M1 ;
        RECT 24.815 17.975 25.065 21.505 ;
  LAYER M1 ;
        RECT 24.815 23.855 25.065 27.385 ;
  LAYER M1 ;
        RECT 24.385 0.335 24.635 3.865 ;
  LAYER M1 ;
        RECT 24.385 4.115 24.635 5.125 ;
  LAYER M1 ;
        RECT 24.385 6.215 24.635 9.745 ;
  LAYER M1 ;
        RECT 24.385 9.995 24.635 11.005 ;
  LAYER M1 ;
        RECT 24.385 12.095 24.635 15.625 ;
  LAYER M1 ;
        RECT 24.385 15.875 24.635 16.885 ;
  LAYER M1 ;
        RECT 24.385 17.975 24.635 21.505 ;
  LAYER M1 ;
        RECT 24.385 21.755 24.635 22.765 ;
  LAYER M1 ;
        RECT 24.385 23.855 24.635 27.385 ;
  LAYER M1 ;
        RECT 24.385 27.635 24.635 28.645 ;
  LAYER M1 ;
        RECT 24.385 29.735 24.635 30.745 ;
  LAYER M1 ;
        RECT 23.955 0.335 24.205 3.865 ;
  LAYER M1 ;
        RECT 23.955 6.215 24.205 9.745 ;
  LAYER M1 ;
        RECT 23.955 12.095 24.205 15.625 ;
  LAYER M1 ;
        RECT 23.955 17.975 24.205 21.505 ;
  LAYER M1 ;
        RECT 23.955 23.855 24.205 27.385 ;
  LAYER M2 ;
        RECT 24.34 0.28 32.42 0.56 ;
  LAYER M2 ;
        RECT 24.34 4.48 32.42 4.76 ;
  LAYER M2 ;
        RECT 23.91 0.7 32.85 0.98 ;
  LAYER M2 ;
        RECT 24.34 6.16 32.42 6.44 ;
  LAYER M2 ;
        RECT 24.34 10.36 32.42 10.64 ;
  LAYER M2 ;
        RECT 23.91 6.58 32.85 6.86 ;
  LAYER M2 ;
        RECT 24.34 12.04 32.42 12.32 ;
  LAYER M2 ;
        RECT 24.34 16.24 32.42 16.52 ;
  LAYER M2 ;
        RECT 23.91 12.46 32.85 12.74 ;
  LAYER M2 ;
        RECT 24.34 17.92 32.42 18.2 ;
  LAYER M2 ;
        RECT 24.34 22.12 32.42 22.4 ;
  LAYER M2 ;
        RECT 23.91 18.34 32.85 18.62 ;
  LAYER M2 ;
        RECT 24.34 23.8 32.42 24.08 ;
  LAYER M2 ;
        RECT 24.34 28 32.42 28.28 ;
  LAYER M2 ;
        RECT 24.34 30.1 32.42 30.38 ;
  LAYER M2 ;
        RECT 23.91 24.22 32.85 24.5 ;
  LAYER M3 ;
        RECT 28.24 0.26 28.52 28.3 ;
  LAYER M3 ;
        RECT 27.81 0.68 28.09 30.4 ;
  LAYER M1 ;
        RECT 1.165 31.415 1.415 34.945 ;
  LAYER M1 ;
        RECT 1.165 35.195 1.415 36.205 ;
  LAYER M1 ;
        RECT 1.165 37.295 1.415 40.825 ;
  LAYER M1 ;
        RECT 1.165 41.075 1.415 42.085 ;
  LAYER M1 ;
        RECT 1.165 43.175 1.415 46.705 ;
  LAYER M1 ;
        RECT 1.165 46.955 1.415 47.965 ;
  LAYER M1 ;
        RECT 1.165 49.055 1.415 52.585 ;
  LAYER M1 ;
        RECT 1.165 52.835 1.415 53.845 ;
  LAYER M1 ;
        RECT 1.165 54.935 1.415 55.945 ;
  LAYER M1 ;
        RECT 0.735 31.415 0.985 34.945 ;
  LAYER M1 ;
        RECT 0.735 37.295 0.985 40.825 ;
  LAYER M1 ;
        RECT 0.735 43.175 0.985 46.705 ;
  LAYER M1 ;
        RECT 0.735 49.055 0.985 52.585 ;
  LAYER M1 ;
        RECT 1.595 31.415 1.845 34.945 ;
  LAYER M1 ;
        RECT 1.595 37.295 1.845 40.825 ;
  LAYER M1 ;
        RECT 1.595 43.175 1.845 46.705 ;
  LAYER M1 ;
        RECT 1.595 49.055 1.845 52.585 ;
  LAYER M1 ;
        RECT 2.025 31.415 2.275 34.945 ;
  LAYER M1 ;
        RECT 2.025 35.195 2.275 36.205 ;
  LAYER M1 ;
        RECT 2.025 37.295 2.275 40.825 ;
  LAYER M1 ;
        RECT 2.025 41.075 2.275 42.085 ;
  LAYER M1 ;
        RECT 2.025 43.175 2.275 46.705 ;
  LAYER M1 ;
        RECT 2.025 46.955 2.275 47.965 ;
  LAYER M1 ;
        RECT 2.025 49.055 2.275 52.585 ;
  LAYER M1 ;
        RECT 2.025 52.835 2.275 53.845 ;
  LAYER M1 ;
        RECT 2.025 54.935 2.275 55.945 ;
  LAYER M1 ;
        RECT 2.455 31.415 2.705 34.945 ;
  LAYER M1 ;
        RECT 2.455 37.295 2.705 40.825 ;
  LAYER M1 ;
        RECT 2.455 43.175 2.705 46.705 ;
  LAYER M1 ;
        RECT 2.455 49.055 2.705 52.585 ;
  LAYER M1 ;
        RECT 2.885 31.415 3.135 34.945 ;
  LAYER M1 ;
        RECT 2.885 35.195 3.135 36.205 ;
  LAYER M1 ;
        RECT 2.885 37.295 3.135 40.825 ;
  LAYER M1 ;
        RECT 2.885 41.075 3.135 42.085 ;
  LAYER M1 ;
        RECT 2.885 43.175 3.135 46.705 ;
  LAYER M1 ;
        RECT 2.885 46.955 3.135 47.965 ;
  LAYER M1 ;
        RECT 2.885 49.055 3.135 52.585 ;
  LAYER M1 ;
        RECT 2.885 52.835 3.135 53.845 ;
  LAYER M1 ;
        RECT 2.885 54.935 3.135 55.945 ;
  LAYER M1 ;
        RECT 3.315 31.415 3.565 34.945 ;
  LAYER M1 ;
        RECT 3.315 37.295 3.565 40.825 ;
  LAYER M1 ;
        RECT 3.315 43.175 3.565 46.705 ;
  LAYER M1 ;
        RECT 3.315 49.055 3.565 52.585 ;
  LAYER M1 ;
        RECT 3.745 31.415 3.995 34.945 ;
  LAYER M1 ;
        RECT 3.745 35.195 3.995 36.205 ;
  LAYER M1 ;
        RECT 3.745 37.295 3.995 40.825 ;
  LAYER M1 ;
        RECT 3.745 41.075 3.995 42.085 ;
  LAYER M1 ;
        RECT 3.745 43.175 3.995 46.705 ;
  LAYER M1 ;
        RECT 3.745 46.955 3.995 47.965 ;
  LAYER M1 ;
        RECT 3.745 49.055 3.995 52.585 ;
  LAYER M1 ;
        RECT 3.745 52.835 3.995 53.845 ;
  LAYER M1 ;
        RECT 3.745 54.935 3.995 55.945 ;
  LAYER M1 ;
        RECT 4.175 31.415 4.425 34.945 ;
  LAYER M1 ;
        RECT 4.175 37.295 4.425 40.825 ;
  LAYER M1 ;
        RECT 4.175 43.175 4.425 46.705 ;
  LAYER M1 ;
        RECT 4.175 49.055 4.425 52.585 ;
  LAYER M1 ;
        RECT 4.605 31.415 4.855 34.945 ;
  LAYER M1 ;
        RECT 4.605 35.195 4.855 36.205 ;
  LAYER M1 ;
        RECT 4.605 37.295 4.855 40.825 ;
  LAYER M1 ;
        RECT 4.605 41.075 4.855 42.085 ;
  LAYER M1 ;
        RECT 4.605 43.175 4.855 46.705 ;
  LAYER M1 ;
        RECT 4.605 46.955 4.855 47.965 ;
  LAYER M1 ;
        RECT 4.605 49.055 4.855 52.585 ;
  LAYER M1 ;
        RECT 4.605 52.835 4.855 53.845 ;
  LAYER M1 ;
        RECT 4.605 54.935 4.855 55.945 ;
  LAYER M1 ;
        RECT 5.035 31.415 5.285 34.945 ;
  LAYER M1 ;
        RECT 5.035 37.295 5.285 40.825 ;
  LAYER M1 ;
        RECT 5.035 43.175 5.285 46.705 ;
  LAYER M1 ;
        RECT 5.035 49.055 5.285 52.585 ;
  LAYER M1 ;
        RECT 5.465 31.415 5.715 34.945 ;
  LAYER M1 ;
        RECT 5.465 35.195 5.715 36.205 ;
  LAYER M1 ;
        RECT 5.465 37.295 5.715 40.825 ;
  LAYER M1 ;
        RECT 5.465 41.075 5.715 42.085 ;
  LAYER M1 ;
        RECT 5.465 43.175 5.715 46.705 ;
  LAYER M1 ;
        RECT 5.465 46.955 5.715 47.965 ;
  LAYER M1 ;
        RECT 5.465 49.055 5.715 52.585 ;
  LAYER M1 ;
        RECT 5.465 52.835 5.715 53.845 ;
  LAYER M1 ;
        RECT 5.465 54.935 5.715 55.945 ;
  LAYER M1 ;
        RECT 5.895 31.415 6.145 34.945 ;
  LAYER M1 ;
        RECT 5.895 37.295 6.145 40.825 ;
  LAYER M1 ;
        RECT 5.895 43.175 6.145 46.705 ;
  LAYER M1 ;
        RECT 5.895 49.055 6.145 52.585 ;
  LAYER M1 ;
        RECT 6.325 31.415 6.575 34.945 ;
  LAYER M1 ;
        RECT 6.325 35.195 6.575 36.205 ;
  LAYER M1 ;
        RECT 6.325 37.295 6.575 40.825 ;
  LAYER M1 ;
        RECT 6.325 41.075 6.575 42.085 ;
  LAYER M1 ;
        RECT 6.325 43.175 6.575 46.705 ;
  LAYER M1 ;
        RECT 6.325 46.955 6.575 47.965 ;
  LAYER M1 ;
        RECT 6.325 49.055 6.575 52.585 ;
  LAYER M1 ;
        RECT 6.325 52.835 6.575 53.845 ;
  LAYER M1 ;
        RECT 6.325 54.935 6.575 55.945 ;
  LAYER M1 ;
        RECT 6.755 31.415 7.005 34.945 ;
  LAYER M1 ;
        RECT 6.755 37.295 7.005 40.825 ;
  LAYER M1 ;
        RECT 6.755 43.175 7.005 46.705 ;
  LAYER M1 ;
        RECT 6.755 49.055 7.005 52.585 ;
  LAYER M1 ;
        RECT 7.185 31.415 7.435 34.945 ;
  LAYER M1 ;
        RECT 7.185 35.195 7.435 36.205 ;
  LAYER M1 ;
        RECT 7.185 37.295 7.435 40.825 ;
  LAYER M1 ;
        RECT 7.185 41.075 7.435 42.085 ;
  LAYER M1 ;
        RECT 7.185 43.175 7.435 46.705 ;
  LAYER M1 ;
        RECT 7.185 46.955 7.435 47.965 ;
  LAYER M1 ;
        RECT 7.185 49.055 7.435 52.585 ;
  LAYER M1 ;
        RECT 7.185 52.835 7.435 53.845 ;
  LAYER M1 ;
        RECT 7.185 54.935 7.435 55.945 ;
  LAYER M1 ;
        RECT 7.615 31.415 7.865 34.945 ;
  LAYER M1 ;
        RECT 7.615 37.295 7.865 40.825 ;
  LAYER M1 ;
        RECT 7.615 43.175 7.865 46.705 ;
  LAYER M1 ;
        RECT 7.615 49.055 7.865 52.585 ;
  LAYER M1 ;
        RECT 8.045 31.415 8.295 34.945 ;
  LAYER M1 ;
        RECT 8.045 35.195 8.295 36.205 ;
  LAYER M1 ;
        RECT 8.045 37.295 8.295 40.825 ;
  LAYER M1 ;
        RECT 8.045 41.075 8.295 42.085 ;
  LAYER M1 ;
        RECT 8.045 43.175 8.295 46.705 ;
  LAYER M1 ;
        RECT 8.045 46.955 8.295 47.965 ;
  LAYER M1 ;
        RECT 8.045 49.055 8.295 52.585 ;
  LAYER M1 ;
        RECT 8.045 52.835 8.295 53.845 ;
  LAYER M1 ;
        RECT 8.045 54.935 8.295 55.945 ;
  LAYER M1 ;
        RECT 8.475 31.415 8.725 34.945 ;
  LAYER M1 ;
        RECT 8.475 37.295 8.725 40.825 ;
  LAYER M1 ;
        RECT 8.475 43.175 8.725 46.705 ;
  LAYER M1 ;
        RECT 8.475 49.055 8.725 52.585 ;
  LAYER M1 ;
        RECT 8.905 31.415 9.155 34.945 ;
  LAYER M1 ;
        RECT 8.905 35.195 9.155 36.205 ;
  LAYER M1 ;
        RECT 8.905 37.295 9.155 40.825 ;
  LAYER M1 ;
        RECT 8.905 41.075 9.155 42.085 ;
  LAYER M1 ;
        RECT 8.905 43.175 9.155 46.705 ;
  LAYER M1 ;
        RECT 8.905 46.955 9.155 47.965 ;
  LAYER M1 ;
        RECT 8.905 49.055 9.155 52.585 ;
  LAYER M1 ;
        RECT 8.905 52.835 9.155 53.845 ;
  LAYER M1 ;
        RECT 8.905 54.935 9.155 55.945 ;
  LAYER M1 ;
        RECT 9.335 31.415 9.585 34.945 ;
  LAYER M1 ;
        RECT 9.335 37.295 9.585 40.825 ;
  LAYER M1 ;
        RECT 9.335 43.175 9.585 46.705 ;
  LAYER M1 ;
        RECT 9.335 49.055 9.585 52.585 ;
  LAYER M1 ;
        RECT 9.765 31.415 10.015 34.945 ;
  LAYER M1 ;
        RECT 9.765 35.195 10.015 36.205 ;
  LAYER M1 ;
        RECT 9.765 37.295 10.015 40.825 ;
  LAYER M1 ;
        RECT 9.765 41.075 10.015 42.085 ;
  LAYER M1 ;
        RECT 9.765 43.175 10.015 46.705 ;
  LAYER M1 ;
        RECT 9.765 46.955 10.015 47.965 ;
  LAYER M1 ;
        RECT 9.765 49.055 10.015 52.585 ;
  LAYER M1 ;
        RECT 9.765 52.835 10.015 53.845 ;
  LAYER M1 ;
        RECT 9.765 54.935 10.015 55.945 ;
  LAYER M1 ;
        RECT 10.195 31.415 10.445 34.945 ;
  LAYER M1 ;
        RECT 10.195 37.295 10.445 40.825 ;
  LAYER M1 ;
        RECT 10.195 43.175 10.445 46.705 ;
  LAYER M1 ;
        RECT 10.195 49.055 10.445 52.585 ;
  LAYER M1 ;
        RECT 10.625 31.415 10.875 34.945 ;
  LAYER M1 ;
        RECT 10.625 35.195 10.875 36.205 ;
  LAYER M1 ;
        RECT 10.625 37.295 10.875 40.825 ;
  LAYER M1 ;
        RECT 10.625 41.075 10.875 42.085 ;
  LAYER M1 ;
        RECT 10.625 43.175 10.875 46.705 ;
  LAYER M1 ;
        RECT 10.625 46.955 10.875 47.965 ;
  LAYER M1 ;
        RECT 10.625 49.055 10.875 52.585 ;
  LAYER M1 ;
        RECT 10.625 52.835 10.875 53.845 ;
  LAYER M1 ;
        RECT 10.625 54.935 10.875 55.945 ;
  LAYER M1 ;
        RECT 11.055 31.415 11.305 34.945 ;
  LAYER M1 ;
        RECT 11.055 37.295 11.305 40.825 ;
  LAYER M1 ;
        RECT 11.055 43.175 11.305 46.705 ;
  LAYER M1 ;
        RECT 11.055 49.055 11.305 52.585 ;
  LAYER M1 ;
        RECT 11.485 31.415 11.735 34.945 ;
  LAYER M1 ;
        RECT 11.485 35.195 11.735 36.205 ;
  LAYER M1 ;
        RECT 11.485 37.295 11.735 40.825 ;
  LAYER M1 ;
        RECT 11.485 41.075 11.735 42.085 ;
  LAYER M1 ;
        RECT 11.485 43.175 11.735 46.705 ;
  LAYER M1 ;
        RECT 11.485 46.955 11.735 47.965 ;
  LAYER M1 ;
        RECT 11.485 49.055 11.735 52.585 ;
  LAYER M1 ;
        RECT 11.485 52.835 11.735 53.845 ;
  LAYER M1 ;
        RECT 11.485 54.935 11.735 55.945 ;
  LAYER M1 ;
        RECT 11.915 31.415 12.165 34.945 ;
  LAYER M1 ;
        RECT 11.915 37.295 12.165 40.825 ;
  LAYER M1 ;
        RECT 11.915 43.175 12.165 46.705 ;
  LAYER M1 ;
        RECT 11.915 49.055 12.165 52.585 ;
  LAYER M1 ;
        RECT 12.345 31.415 12.595 34.945 ;
  LAYER M1 ;
        RECT 12.345 35.195 12.595 36.205 ;
  LAYER M1 ;
        RECT 12.345 37.295 12.595 40.825 ;
  LAYER M1 ;
        RECT 12.345 41.075 12.595 42.085 ;
  LAYER M1 ;
        RECT 12.345 43.175 12.595 46.705 ;
  LAYER M1 ;
        RECT 12.345 46.955 12.595 47.965 ;
  LAYER M1 ;
        RECT 12.345 49.055 12.595 52.585 ;
  LAYER M1 ;
        RECT 12.345 52.835 12.595 53.845 ;
  LAYER M1 ;
        RECT 12.345 54.935 12.595 55.945 ;
  LAYER M1 ;
        RECT 12.775 31.415 13.025 34.945 ;
  LAYER M1 ;
        RECT 12.775 37.295 13.025 40.825 ;
  LAYER M1 ;
        RECT 12.775 43.175 13.025 46.705 ;
  LAYER M1 ;
        RECT 12.775 49.055 13.025 52.585 ;
  LAYER M1 ;
        RECT 13.205 31.415 13.455 34.945 ;
  LAYER M1 ;
        RECT 13.205 35.195 13.455 36.205 ;
  LAYER M1 ;
        RECT 13.205 37.295 13.455 40.825 ;
  LAYER M1 ;
        RECT 13.205 41.075 13.455 42.085 ;
  LAYER M1 ;
        RECT 13.205 43.175 13.455 46.705 ;
  LAYER M1 ;
        RECT 13.205 46.955 13.455 47.965 ;
  LAYER M1 ;
        RECT 13.205 49.055 13.455 52.585 ;
  LAYER M1 ;
        RECT 13.205 52.835 13.455 53.845 ;
  LAYER M1 ;
        RECT 13.205 54.935 13.455 55.945 ;
  LAYER M1 ;
        RECT 13.635 31.415 13.885 34.945 ;
  LAYER M1 ;
        RECT 13.635 37.295 13.885 40.825 ;
  LAYER M1 ;
        RECT 13.635 43.175 13.885 46.705 ;
  LAYER M1 ;
        RECT 13.635 49.055 13.885 52.585 ;
  LAYER M1 ;
        RECT 14.065 31.415 14.315 34.945 ;
  LAYER M1 ;
        RECT 14.065 35.195 14.315 36.205 ;
  LAYER M1 ;
        RECT 14.065 37.295 14.315 40.825 ;
  LAYER M1 ;
        RECT 14.065 41.075 14.315 42.085 ;
  LAYER M1 ;
        RECT 14.065 43.175 14.315 46.705 ;
  LAYER M1 ;
        RECT 14.065 46.955 14.315 47.965 ;
  LAYER M1 ;
        RECT 14.065 49.055 14.315 52.585 ;
  LAYER M1 ;
        RECT 14.065 52.835 14.315 53.845 ;
  LAYER M1 ;
        RECT 14.065 54.935 14.315 55.945 ;
  LAYER M1 ;
        RECT 14.495 31.415 14.745 34.945 ;
  LAYER M1 ;
        RECT 14.495 37.295 14.745 40.825 ;
  LAYER M1 ;
        RECT 14.495 43.175 14.745 46.705 ;
  LAYER M1 ;
        RECT 14.495 49.055 14.745 52.585 ;
  LAYER M1 ;
        RECT 14.925 31.415 15.175 34.945 ;
  LAYER M1 ;
        RECT 14.925 35.195 15.175 36.205 ;
  LAYER M1 ;
        RECT 14.925 37.295 15.175 40.825 ;
  LAYER M1 ;
        RECT 14.925 41.075 15.175 42.085 ;
  LAYER M1 ;
        RECT 14.925 43.175 15.175 46.705 ;
  LAYER M1 ;
        RECT 14.925 46.955 15.175 47.965 ;
  LAYER M1 ;
        RECT 14.925 49.055 15.175 52.585 ;
  LAYER M1 ;
        RECT 14.925 52.835 15.175 53.845 ;
  LAYER M1 ;
        RECT 14.925 54.935 15.175 55.945 ;
  LAYER M1 ;
        RECT 15.355 31.415 15.605 34.945 ;
  LAYER M1 ;
        RECT 15.355 37.295 15.605 40.825 ;
  LAYER M1 ;
        RECT 15.355 43.175 15.605 46.705 ;
  LAYER M1 ;
        RECT 15.355 49.055 15.605 52.585 ;
  LAYER M1 ;
        RECT 15.785 31.415 16.035 34.945 ;
  LAYER M1 ;
        RECT 15.785 35.195 16.035 36.205 ;
  LAYER M1 ;
        RECT 15.785 37.295 16.035 40.825 ;
  LAYER M1 ;
        RECT 15.785 41.075 16.035 42.085 ;
  LAYER M1 ;
        RECT 15.785 43.175 16.035 46.705 ;
  LAYER M1 ;
        RECT 15.785 46.955 16.035 47.965 ;
  LAYER M1 ;
        RECT 15.785 49.055 16.035 52.585 ;
  LAYER M1 ;
        RECT 15.785 52.835 16.035 53.845 ;
  LAYER M1 ;
        RECT 15.785 54.935 16.035 55.945 ;
  LAYER M1 ;
        RECT 16.215 31.415 16.465 34.945 ;
  LAYER M1 ;
        RECT 16.215 37.295 16.465 40.825 ;
  LAYER M1 ;
        RECT 16.215 43.175 16.465 46.705 ;
  LAYER M1 ;
        RECT 16.215 49.055 16.465 52.585 ;
  LAYER M1 ;
        RECT 16.645 31.415 16.895 34.945 ;
  LAYER M1 ;
        RECT 16.645 35.195 16.895 36.205 ;
  LAYER M1 ;
        RECT 16.645 37.295 16.895 40.825 ;
  LAYER M1 ;
        RECT 16.645 41.075 16.895 42.085 ;
  LAYER M1 ;
        RECT 16.645 43.175 16.895 46.705 ;
  LAYER M1 ;
        RECT 16.645 46.955 16.895 47.965 ;
  LAYER M1 ;
        RECT 16.645 49.055 16.895 52.585 ;
  LAYER M1 ;
        RECT 16.645 52.835 16.895 53.845 ;
  LAYER M1 ;
        RECT 16.645 54.935 16.895 55.945 ;
  LAYER M1 ;
        RECT 17.075 31.415 17.325 34.945 ;
  LAYER M1 ;
        RECT 17.075 37.295 17.325 40.825 ;
  LAYER M1 ;
        RECT 17.075 43.175 17.325 46.705 ;
  LAYER M1 ;
        RECT 17.075 49.055 17.325 52.585 ;
  LAYER M1 ;
        RECT 17.505 31.415 17.755 34.945 ;
  LAYER M1 ;
        RECT 17.505 35.195 17.755 36.205 ;
  LAYER M1 ;
        RECT 17.505 37.295 17.755 40.825 ;
  LAYER M1 ;
        RECT 17.505 41.075 17.755 42.085 ;
  LAYER M1 ;
        RECT 17.505 43.175 17.755 46.705 ;
  LAYER M1 ;
        RECT 17.505 46.955 17.755 47.965 ;
  LAYER M1 ;
        RECT 17.505 49.055 17.755 52.585 ;
  LAYER M1 ;
        RECT 17.505 52.835 17.755 53.845 ;
  LAYER M1 ;
        RECT 17.505 54.935 17.755 55.945 ;
  LAYER M1 ;
        RECT 17.935 31.415 18.185 34.945 ;
  LAYER M1 ;
        RECT 17.935 37.295 18.185 40.825 ;
  LAYER M1 ;
        RECT 17.935 43.175 18.185 46.705 ;
  LAYER M1 ;
        RECT 17.935 49.055 18.185 52.585 ;
  LAYER M1 ;
        RECT 18.365 31.415 18.615 34.945 ;
  LAYER M1 ;
        RECT 18.365 35.195 18.615 36.205 ;
  LAYER M1 ;
        RECT 18.365 37.295 18.615 40.825 ;
  LAYER M1 ;
        RECT 18.365 41.075 18.615 42.085 ;
  LAYER M1 ;
        RECT 18.365 43.175 18.615 46.705 ;
  LAYER M1 ;
        RECT 18.365 46.955 18.615 47.965 ;
  LAYER M1 ;
        RECT 18.365 49.055 18.615 52.585 ;
  LAYER M1 ;
        RECT 18.365 52.835 18.615 53.845 ;
  LAYER M1 ;
        RECT 18.365 54.935 18.615 55.945 ;
  LAYER M1 ;
        RECT 18.795 31.415 19.045 34.945 ;
  LAYER M1 ;
        RECT 18.795 37.295 19.045 40.825 ;
  LAYER M1 ;
        RECT 18.795 43.175 19.045 46.705 ;
  LAYER M1 ;
        RECT 18.795 49.055 19.045 52.585 ;
  LAYER M1 ;
        RECT 19.225 31.415 19.475 34.945 ;
  LAYER M1 ;
        RECT 19.225 35.195 19.475 36.205 ;
  LAYER M1 ;
        RECT 19.225 37.295 19.475 40.825 ;
  LAYER M1 ;
        RECT 19.225 41.075 19.475 42.085 ;
  LAYER M1 ;
        RECT 19.225 43.175 19.475 46.705 ;
  LAYER M1 ;
        RECT 19.225 46.955 19.475 47.965 ;
  LAYER M1 ;
        RECT 19.225 49.055 19.475 52.585 ;
  LAYER M1 ;
        RECT 19.225 52.835 19.475 53.845 ;
  LAYER M1 ;
        RECT 19.225 54.935 19.475 55.945 ;
  LAYER M1 ;
        RECT 19.655 31.415 19.905 34.945 ;
  LAYER M1 ;
        RECT 19.655 37.295 19.905 40.825 ;
  LAYER M1 ;
        RECT 19.655 43.175 19.905 46.705 ;
  LAYER M1 ;
        RECT 19.655 49.055 19.905 52.585 ;
  LAYER M1 ;
        RECT 20.085 31.415 20.335 34.945 ;
  LAYER M1 ;
        RECT 20.085 35.195 20.335 36.205 ;
  LAYER M1 ;
        RECT 20.085 37.295 20.335 40.825 ;
  LAYER M1 ;
        RECT 20.085 41.075 20.335 42.085 ;
  LAYER M1 ;
        RECT 20.085 43.175 20.335 46.705 ;
  LAYER M1 ;
        RECT 20.085 46.955 20.335 47.965 ;
  LAYER M1 ;
        RECT 20.085 49.055 20.335 52.585 ;
  LAYER M1 ;
        RECT 20.085 52.835 20.335 53.845 ;
  LAYER M1 ;
        RECT 20.085 54.935 20.335 55.945 ;
  LAYER M1 ;
        RECT 20.515 31.415 20.765 34.945 ;
  LAYER M1 ;
        RECT 20.515 37.295 20.765 40.825 ;
  LAYER M1 ;
        RECT 20.515 43.175 20.765 46.705 ;
  LAYER M1 ;
        RECT 20.515 49.055 20.765 52.585 ;
  LAYER M1 ;
        RECT 20.945 31.415 21.195 34.945 ;
  LAYER M1 ;
        RECT 20.945 35.195 21.195 36.205 ;
  LAYER M1 ;
        RECT 20.945 37.295 21.195 40.825 ;
  LAYER M1 ;
        RECT 20.945 41.075 21.195 42.085 ;
  LAYER M1 ;
        RECT 20.945 43.175 21.195 46.705 ;
  LAYER M1 ;
        RECT 20.945 46.955 21.195 47.965 ;
  LAYER M1 ;
        RECT 20.945 49.055 21.195 52.585 ;
  LAYER M1 ;
        RECT 20.945 52.835 21.195 53.845 ;
  LAYER M1 ;
        RECT 20.945 54.935 21.195 55.945 ;
  LAYER M1 ;
        RECT 21.375 31.415 21.625 34.945 ;
  LAYER M1 ;
        RECT 21.375 37.295 21.625 40.825 ;
  LAYER M1 ;
        RECT 21.375 43.175 21.625 46.705 ;
  LAYER M1 ;
        RECT 21.375 49.055 21.625 52.585 ;
  LAYER M1 ;
        RECT 21.805 31.415 22.055 34.945 ;
  LAYER M1 ;
        RECT 21.805 35.195 22.055 36.205 ;
  LAYER M1 ;
        RECT 21.805 37.295 22.055 40.825 ;
  LAYER M1 ;
        RECT 21.805 41.075 22.055 42.085 ;
  LAYER M1 ;
        RECT 21.805 43.175 22.055 46.705 ;
  LAYER M1 ;
        RECT 21.805 46.955 22.055 47.965 ;
  LAYER M1 ;
        RECT 21.805 49.055 22.055 52.585 ;
  LAYER M1 ;
        RECT 21.805 52.835 22.055 53.845 ;
  LAYER M1 ;
        RECT 21.805 54.935 22.055 55.945 ;
  LAYER M1 ;
        RECT 22.235 31.415 22.485 34.945 ;
  LAYER M1 ;
        RECT 22.235 37.295 22.485 40.825 ;
  LAYER M1 ;
        RECT 22.235 43.175 22.485 46.705 ;
  LAYER M1 ;
        RECT 22.235 49.055 22.485 52.585 ;
  LAYER M1 ;
        RECT 22.665 31.415 22.915 34.945 ;
  LAYER M1 ;
        RECT 22.665 35.195 22.915 36.205 ;
  LAYER M1 ;
        RECT 22.665 37.295 22.915 40.825 ;
  LAYER M1 ;
        RECT 22.665 41.075 22.915 42.085 ;
  LAYER M1 ;
        RECT 22.665 43.175 22.915 46.705 ;
  LAYER M1 ;
        RECT 22.665 46.955 22.915 47.965 ;
  LAYER M1 ;
        RECT 22.665 49.055 22.915 52.585 ;
  LAYER M1 ;
        RECT 22.665 52.835 22.915 53.845 ;
  LAYER M1 ;
        RECT 22.665 54.935 22.915 55.945 ;
  LAYER M1 ;
        RECT 23.095 31.415 23.345 34.945 ;
  LAYER M1 ;
        RECT 23.095 37.295 23.345 40.825 ;
  LAYER M1 ;
        RECT 23.095 43.175 23.345 46.705 ;
  LAYER M1 ;
        RECT 23.095 49.055 23.345 52.585 ;
  LAYER M1 ;
        RECT 23.525 31.415 23.775 34.945 ;
  LAYER M1 ;
        RECT 23.525 35.195 23.775 36.205 ;
  LAYER M1 ;
        RECT 23.525 37.295 23.775 40.825 ;
  LAYER M1 ;
        RECT 23.525 41.075 23.775 42.085 ;
  LAYER M1 ;
        RECT 23.525 43.175 23.775 46.705 ;
  LAYER M1 ;
        RECT 23.525 46.955 23.775 47.965 ;
  LAYER M1 ;
        RECT 23.525 49.055 23.775 52.585 ;
  LAYER M1 ;
        RECT 23.525 52.835 23.775 53.845 ;
  LAYER M1 ;
        RECT 23.525 54.935 23.775 55.945 ;
  LAYER M1 ;
        RECT 23.955 31.415 24.205 34.945 ;
  LAYER M1 ;
        RECT 23.955 37.295 24.205 40.825 ;
  LAYER M1 ;
        RECT 23.955 43.175 24.205 46.705 ;
  LAYER M1 ;
        RECT 23.955 49.055 24.205 52.585 ;
  LAYER M1 ;
        RECT 24.385 31.415 24.635 34.945 ;
  LAYER M1 ;
        RECT 24.385 35.195 24.635 36.205 ;
  LAYER M1 ;
        RECT 24.385 37.295 24.635 40.825 ;
  LAYER M1 ;
        RECT 24.385 41.075 24.635 42.085 ;
  LAYER M1 ;
        RECT 24.385 43.175 24.635 46.705 ;
  LAYER M1 ;
        RECT 24.385 46.955 24.635 47.965 ;
  LAYER M1 ;
        RECT 24.385 49.055 24.635 52.585 ;
  LAYER M1 ;
        RECT 24.385 52.835 24.635 53.845 ;
  LAYER M1 ;
        RECT 24.385 54.935 24.635 55.945 ;
  LAYER M1 ;
        RECT 24.815 31.415 25.065 34.945 ;
  LAYER M1 ;
        RECT 24.815 37.295 25.065 40.825 ;
  LAYER M1 ;
        RECT 24.815 43.175 25.065 46.705 ;
  LAYER M1 ;
        RECT 24.815 49.055 25.065 52.585 ;
  LAYER M1 ;
        RECT 25.245 31.415 25.495 34.945 ;
  LAYER M1 ;
        RECT 25.245 35.195 25.495 36.205 ;
  LAYER M1 ;
        RECT 25.245 37.295 25.495 40.825 ;
  LAYER M1 ;
        RECT 25.245 41.075 25.495 42.085 ;
  LAYER M1 ;
        RECT 25.245 43.175 25.495 46.705 ;
  LAYER M1 ;
        RECT 25.245 46.955 25.495 47.965 ;
  LAYER M1 ;
        RECT 25.245 49.055 25.495 52.585 ;
  LAYER M1 ;
        RECT 25.245 52.835 25.495 53.845 ;
  LAYER M1 ;
        RECT 25.245 54.935 25.495 55.945 ;
  LAYER M1 ;
        RECT 25.675 31.415 25.925 34.945 ;
  LAYER M1 ;
        RECT 25.675 37.295 25.925 40.825 ;
  LAYER M1 ;
        RECT 25.675 43.175 25.925 46.705 ;
  LAYER M1 ;
        RECT 25.675 49.055 25.925 52.585 ;
  LAYER M1 ;
        RECT 26.105 31.415 26.355 34.945 ;
  LAYER M1 ;
        RECT 26.105 35.195 26.355 36.205 ;
  LAYER M1 ;
        RECT 26.105 37.295 26.355 40.825 ;
  LAYER M1 ;
        RECT 26.105 41.075 26.355 42.085 ;
  LAYER M1 ;
        RECT 26.105 43.175 26.355 46.705 ;
  LAYER M1 ;
        RECT 26.105 46.955 26.355 47.965 ;
  LAYER M1 ;
        RECT 26.105 49.055 26.355 52.585 ;
  LAYER M1 ;
        RECT 26.105 52.835 26.355 53.845 ;
  LAYER M1 ;
        RECT 26.105 54.935 26.355 55.945 ;
  LAYER M1 ;
        RECT 26.535 31.415 26.785 34.945 ;
  LAYER M1 ;
        RECT 26.535 37.295 26.785 40.825 ;
  LAYER M1 ;
        RECT 26.535 43.175 26.785 46.705 ;
  LAYER M1 ;
        RECT 26.535 49.055 26.785 52.585 ;
  LAYER M1 ;
        RECT 26.965 31.415 27.215 34.945 ;
  LAYER M1 ;
        RECT 26.965 35.195 27.215 36.205 ;
  LAYER M1 ;
        RECT 26.965 37.295 27.215 40.825 ;
  LAYER M1 ;
        RECT 26.965 41.075 27.215 42.085 ;
  LAYER M1 ;
        RECT 26.965 43.175 27.215 46.705 ;
  LAYER M1 ;
        RECT 26.965 46.955 27.215 47.965 ;
  LAYER M1 ;
        RECT 26.965 49.055 27.215 52.585 ;
  LAYER M1 ;
        RECT 26.965 52.835 27.215 53.845 ;
  LAYER M1 ;
        RECT 26.965 54.935 27.215 55.945 ;
  LAYER M1 ;
        RECT 27.395 31.415 27.645 34.945 ;
  LAYER M1 ;
        RECT 27.395 37.295 27.645 40.825 ;
  LAYER M1 ;
        RECT 27.395 43.175 27.645 46.705 ;
  LAYER M1 ;
        RECT 27.395 49.055 27.645 52.585 ;
  LAYER M1 ;
        RECT 27.825 31.415 28.075 34.945 ;
  LAYER M1 ;
        RECT 27.825 35.195 28.075 36.205 ;
  LAYER M1 ;
        RECT 27.825 37.295 28.075 40.825 ;
  LAYER M1 ;
        RECT 27.825 41.075 28.075 42.085 ;
  LAYER M1 ;
        RECT 27.825 43.175 28.075 46.705 ;
  LAYER M1 ;
        RECT 27.825 46.955 28.075 47.965 ;
  LAYER M1 ;
        RECT 27.825 49.055 28.075 52.585 ;
  LAYER M1 ;
        RECT 27.825 52.835 28.075 53.845 ;
  LAYER M1 ;
        RECT 27.825 54.935 28.075 55.945 ;
  LAYER M1 ;
        RECT 28.255 31.415 28.505 34.945 ;
  LAYER M1 ;
        RECT 28.255 37.295 28.505 40.825 ;
  LAYER M1 ;
        RECT 28.255 43.175 28.505 46.705 ;
  LAYER M1 ;
        RECT 28.255 49.055 28.505 52.585 ;
  LAYER M1 ;
        RECT 28.685 31.415 28.935 34.945 ;
  LAYER M1 ;
        RECT 28.685 35.195 28.935 36.205 ;
  LAYER M1 ;
        RECT 28.685 37.295 28.935 40.825 ;
  LAYER M1 ;
        RECT 28.685 41.075 28.935 42.085 ;
  LAYER M1 ;
        RECT 28.685 43.175 28.935 46.705 ;
  LAYER M1 ;
        RECT 28.685 46.955 28.935 47.965 ;
  LAYER M1 ;
        RECT 28.685 49.055 28.935 52.585 ;
  LAYER M1 ;
        RECT 28.685 52.835 28.935 53.845 ;
  LAYER M1 ;
        RECT 28.685 54.935 28.935 55.945 ;
  LAYER M1 ;
        RECT 29.115 31.415 29.365 34.945 ;
  LAYER M1 ;
        RECT 29.115 37.295 29.365 40.825 ;
  LAYER M1 ;
        RECT 29.115 43.175 29.365 46.705 ;
  LAYER M1 ;
        RECT 29.115 49.055 29.365 52.585 ;
  LAYER M1 ;
        RECT 29.545 31.415 29.795 34.945 ;
  LAYER M1 ;
        RECT 29.545 35.195 29.795 36.205 ;
  LAYER M1 ;
        RECT 29.545 37.295 29.795 40.825 ;
  LAYER M1 ;
        RECT 29.545 41.075 29.795 42.085 ;
  LAYER M1 ;
        RECT 29.545 43.175 29.795 46.705 ;
  LAYER M1 ;
        RECT 29.545 46.955 29.795 47.965 ;
  LAYER M1 ;
        RECT 29.545 49.055 29.795 52.585 ;
  LAYER M1 ;
        RECT 29.545 52.835 29.795 53.845 ;
  LAYER M1 ;
        RECT 29.545 54.935 29.795 55.945 ;
  LAYER M1 ;
        RECT 29.975 31.415 30.225 34.945 ;
  LAYER M1 ;
        RECT 29.975 37.295 30.225 40.825 ;
  LAYER M1 ;
        RECT 29.975 43.175 30.225 46.705 ;
  LAYER M1 ;
        RECT 29.975 49.055 30.225 52.585 ;
  LAYER M1 ;
        RECT 30.405 31.415 30.655 34.945 ;
  LAYER M1 ;
        RECT 30.405 35.195 30.655 36.205 ;
  LAYER M1 ;
        RECT 30.405 37.295 30.655 40.825 ;
  LAYER M1 ;
        RECT 30.405 41.075 30.655 42.085 ;
  LAYER M1 ;
        RECT 30.405 43.175 30.655 46.705 ;
  LAYER M1 ;
        RECT 30.405 46.955 30.655 47.965 ;
  LAYER M1 ;
        RECT 30.405 49.055 30.655 52.585 ;
  LAYER M1 ;
        RECT 30.405 52.835 30.655 53.845 ;
  LAYER M1 ;
        RECT 30.405 54.935 30.655 55.945 ;
  LAYER M1 ;
        RECT 30.835 31.415 31.085 34.945 ;
  LAYER M1 ;
        RECT 30.835 37.295 31.085 40.825 ;
  LAYER M1 ;
        RECT 30.835 43.175 31.085 46.705 ;
  LAYER M1 ;
        RECT 30.835 49.055 31.085 52.585 ;
  LAYER M1 ;
        RECT 31.265 31.415 31.515 34.945 ;
  LAYER M1 ;
        RECT 31.265 35.195 31.515 36.205 ;
  LAYER M1 ;
        RECT 31.265 37.295 31.515 40.825 ;
  LAYER M1 ;
        RECT 31.265 41.075 31.515 42.085 ;
  LAYER M1 ;
        RECT 31.265 43.175 31.515 46.705 ;
  LAYER M1 ;
        RECT 31.265 46.955 31.515 47.965 ;
  LAYER M1 ;
        RECT 31.265 49.055 31.515 52.585 ;
  LAYER M1 ;
        RECT 31.265 52.835 31.515 53.845 ;
  LAYER M1 ;
        RECT 31.265 54.935 31.515 55.945 ;
  LAYER M1 ;
        RECT 31.695 31.415 31.945 34.945 ;
  LAYER M1 ;
        RECT 31.695 37.295 31.945 40.825 ;
  LAYER M1 ;
        RECT 31.695 43.175 31.945 46.705 ;
  LAYER M1 ;
        RECT 31.695 49.055 31.945 52.585 ;
  LAYER M1 ;
        RECT 32.125 31.415 32.375 34.945 ;
  LAYER M1 ;
        RECT 32.125 35.195 32.375 36.205 ;
  LAYER M1 ;
        RECT 32.125 37.295 32.375 40.825 ;
  LAYER M1 ;
        RECT 32.125 41.075 32.375 42.085 ;
  LAYER M1 ;
        RECT 32.125 43.175 32.375 46.705 ;
  LAYER M1 ;
        RECT 32.125 46.955 32.375 47.965 ;
  LAYER M1 ;
        RECT 32.125 49.055 32.375 52.585 ;
  LAYER M1 ;
        RECT 32.125 52.835 32.375 53.845 ;
  LAYER M1 ;
        RECT 32.125 54.935 32.375 55.945 ;
  LAYER M1 ;
        RECT 32.555 31.415 32.805 34.945 ;
  LAYER M1 ;
        RECT 32.555 37.295 32.805 40.825 ;
  LAYER M1 ;
        RECT 32.555 43.175 32.805 46.705 ;
  LAYER M1 ;
        RECT 32.555 49.055 32.805 52.585 ;
  LAYER M2 ;
        RECT 1.12 31.36 32.42 31.64 ;
  LAYER M2 ;
        RECT 1.12 35.56 32.42 35.84 ;
  LAYER M2 ;
        RECT 0.69 31.78 32.85 32.06 ;
  LAYER M2 ;
        RECT 1.12 37.24 32.42 37.52 ;
  LAYER M2 ;
        RECT 1.12 41.44 32.42 41.72 ;
  LAYER M2 ;
        RECT 0.69 37.66 32.85 37.94 ;
  LAYER M2 ;
        RECT 1.12 43.12 32.42 43.4 ;
  LAYER M2 ;
        RECT 1.12 47.32 32.42 47.6 ;
  LAYER M2 ;
        RECT 0.69 43.54 32.85 43.82 ;
  LAYER M2 ;
        RECT 1.12 49 32.42 49.28 ;
  LAYER M2 ;
        RECT 1.12 53.2 32.42 53.48 ;
  LAYER M2 ;
        RECT 1.12 55.3 32.42 55.58 ;
  LAYER M2 ;
        RECT 0.69 49.42 32.85 49.7 ;
  LAYER M3 ;
        RECT 16.63 31.34 16.91 53.5 ;
  LAYER M3 ;
        RECT 17.06 31.76 17.34 55.6 ;
  LAYER M1 ;
        RECT 2.885 16.295 3.135 19.825 ;
  LAYER M1 ;
        RECT 2.885 20.075 3.135 21.085 ;
  LAYER M1 ;
        RECT 2.885 22.175 3.135 25.705 ;
  LAYER M1 ;
        RECT 2.885 25.955 3.135 26.965 ;
  LAYER M1 ;
        RECT 2.885 28.055 3.135 29.065 ;
  LAYER M1 ;
        RECT 3.315 16.295 3.565 19.825 ;
  LAYER M1 ;
        RECT 3.315 22.175 3.565 25.705 ;
  LAYER M1 ;
        RECT 2.455 16.295 2.705 19.825 ;
  LAYER M1 ;
        RECT 2.455 22.175 2.705 25.705 ;
  LAYER M1 ;
        RECT 2.025 16.295 2.275 19.825 ;
  LAYER M1 ;
        RECT 2.025 20.075 2.275 21.085 ;
  LAYER M1 ;
        RECT 2.025 22.175 2.275 25.705 ;
  LAYER M1 ;
        RECT 2.025 25.955 2.275 26.965 ;
  LAYER M1 ;
        RECT 2.025 28.055 2.275 29.065 ;
  LAYER M1 ;
        RECT 1.595 16.295 1.845 19.825 ;
  LAYER M1 ;
        RECT 1.595 22.175 1.845 25.705 ;
  LAYER M1 ;
        RECT 1.165 16.295 1.415 19.825 ;
  LAYER M1 ;
        RECT 1.165 20.075 1.415 21.085 ;
  LAYER M1 ;
        RECT 1.165 22.175 1.415 25.705 ;
  LAYER M1 ;
        RECT 1.165 25.955 1.415 26.965 ;
  LAYER M1 ;
        RECT 1.165 28.055 1.415 29.065 ;
  LAYER M1 ;
        RECT 0.735 16.295 0.985 19.825 ;
  LAYER M1 ;
        RECT 0.735 22.175 0.985 25.705 ;
  LAYER M2 ;
        RECT 1.12 16.24 3.18 16.52 ;
  LAYER M2 ;
        RECT 1.12 20.44 3.18 20.72 ;
  LAYER M2 ;
        RECT 0.69 16.66 3.61 16.94 ;
  LAYER M2 ;
        RECT 1.12 22.12 3.18 22.4 ;
  LAYER M2 ;
        RECT 1.12 26.32 3.18 26.6 ;
  LAYER M2 ;
        RECT 1.12 28.42 3.18 28.7 ;
  LAYER M2 ;
        RECT 0.69 22.54 3.61 22.82 ;
  LAYER M3 ;
        RECT 2.01 16.22 2.29 26.62 ;
  LAYER M3 ;
        RECT 1.58 16.64 1.86 28.72 ;
  LAYER M1 ;
        RECT 63.945 16.295 64.195 19.825 ;
  LAYER M1 ;
        RECT 63.945 20.075 64.195 21.085 ;
  LAYER M1 ;
        RECT 63.945 22.175 64.195 25.705 ;
  LAYER M1 ;
        RECT 63.945 25.955 64.195 26.965 ;
  LAYER M1 ;
        RECT 63.945 28.055 64.195 29.065 ;
  LAYER M1 ;
        RECT 63.515 16.295 63.765 19.825 ;
  LAYER M1 ;
        RECT 63.515 22.175 63.765 25.705 ;
  LAYER M1 ;
        RECT 64.375 16.295 64.625 19.825 ;
  LAYER M1 ;
        RECT 64.375 22.175 64.625 25.705 ;
  LAYER M1 ;
        RECT 64.805 16.295 65.055 19.825 ;
  LAYER M1 ;
        RECT 64.805 20.075 65.055 21.085 ;
  LAYER M1 ;
        RECT 64.805 22.175 65.055 25.705 ;
  LAYER M1 ;
        RECT 64.805 25.955 65.055 26.965 ;
  LAYER M1 ;
        RECT 64.805 28.055 65.055 29.065 ;
  LAYER M1 ;
        RECT 65.235 16.295 65.485 19.825 ;
  LAYER M1 ;
        RECT 65.235 22.175 65.485 25.705 ;
  LAYER M1 ;
        RECT 65.665 16.295 65.915 19.825 ;
  LAYER M1 ;
        RECT 65.665 20.075 65.915 21.085 ;
  LAYER M1 ;
        RECT 65.665 22.175 65.915 25.705 ;
  LAYER M1 ;
        RECT 65.665 25.955 65.915 26.965 ;
  LAYER M1 ;
        RECT 65.665 28.055 65.915 29.065 ;
  LAYER M1 ;
        RECT 66.095 16.295 66.345 19.825 ;
  LAYER M1 ;
        RECT 66.095 22.175 66.345 25.705 ;
  LAYER M2 ;
        RECT 63.9 16.24 65.96 16.52 ;
  LAYER M2 ;
        RECT 63.9 20.44 65.96 20.72 ;
  LAYER M2 ;
        RECT 63.47 16.66 66.39 16.94 ;
  LAYER M2 ;
        RECT 63.9 22.12 65.96 22.4 ;
  LAYER M2 ;
        RECT 63.9 26.32 65.96 26.6 ;
  LAYER M2 ;
        RECT 63.9 28.42 65.96 28.7 ;
  LAYER M2 ;
        RECT 63.47 22.54 66.39 22.82 ;
  LAYER M3 ;
        RECT 64.79 16.22 65.07 26.62 ;
  LAYER M3 ;
        RECT 65.22 16.64 65.5 28.72 ;
  LAYER M1 ;
        RECT 65.665 31.415 65.915 34.945 ;
  LAYER M1 ;
        RECT 65.665 35.195 65.915 36.205 ;
  LAYER M1 ;
        RECT 65.665 37.295 65.915 40.825 ;
  LAYER M1 ;
        RECT 65.665 41.075 65.915 42.085 ;
  LAYER M1 ;
        RECT 65.665 43.175 65.915 46.705 ;
  LAYER M1 ;
        RECT 65.665 46.955 65.915 47.965 ;
  LAYER M1 ;
        RECT 65.665 49.055 65.915 52.585 ;
  LAYER M1 ;
        RECT 65.665 52.835 65.915 53.845 ;
  LAYER M1 ;
        RECT 65.665 54.935 65.915 55.945 ;
  LAYER M1 ;
        RECT 66.095 31.415 66.345 34.945 ;
  LAYER M1 ;
        RECT 66.095 37.295 66.345 40.825 ;
  LAYER M1 ;
        RECT 66.095 43.175 66.345 46.705 ;
  LAYER M1 ;
        RECT 66.095 49.055 66.345 52.585 ;
  LAYER M1 ;
        RECT 65.235 31.415 65.485 34.945 ;
  LAYER M1 ;
        RECT 65.235 37.295 65.485 40.825 ;
  LAYER M1 ;
        RECT 65.235 43.175 65.485 46.705 ;
  LAYER M1 ;
        RECT 65.235 49.055 65.485 52.585 ;
  LAYER M1 ;
        RECT 64.805 31.415 65.055 34.945 ;
  LAYER M1 ;
        RECT 64.805 35.195 65.055 36.205 ;
  LAYER M1 ;
        RECT 64.805 37.295 65.055 40.825 ;
  LAYER M1 ;
        RECT 64.805 41.075 65.055 42.085 ;
  LAYER M1 ;
        RECT 64.805 43.175 65.055 46.705 ;
  LAYER M1 ;
        RECT 64.805 46.955 65.055 47.965 ;
  LAYER M1 ;
        RECT 64.805 49.055 65.055 52.585 ;
  LAYER M1 ;
        RECT 64.805 52.835 65.055 53.845 ;
  LAYER M1 ;
        RECT 64.805 54.935 65.055 55.945 ;
  LAYER M1 ;
        RECT 64.375 31.415 64.625 34.945 ;
  LAYER M1 ;
        RECT 64.375 37.295 64.625 40.825 ;
  LAYER M1 ;
        RECT 64.375 43.175 64.625 46.705 ;
  LAYER M1 ;
        RECT 64.375 49.055 64.625 52.585 ;
  LAYER M1 ;
        RECT 63.945 31.415 64.195 34.945 ;
  LAYER M1 ;
        RECT 63.945 35.195 64.195 36.205 ;
  LAYER M1 ;
        RECT 63.945 37.295 64.195 40.825 ;
  LAYER M1 ;
        RECT 63.945 41.075 64.195 42.085 ;
  LAYER M1 ;
        RECT 63.945 43.175 64.195 46.705 ;
  LAYER M1 ;
        RECT 63.945 46.955 64.195 47.965 ;
  LAYER M1 ;
        RECT 63.945 49.055 64.195 52.585 ;
  LAYER M1 ;
        RECT 63.945 52.835 64.195 53.845 ;
  LAYER M1 ;
        RECT 63.945 54.935 64.195 55.945 ;
  LAYER M1 ;
        RECT 63.515 31.415 63.765 34.945 ;
  LAYER M1 ;
        RECT 63.515 37.295 63.765 40.825 ;
  LAYER M1 ;
        RECT 63.515 43.175 63.765 46.705 ;
  LAYER M1 ;
        RECT 63.515 49.055 63.765 52.585 ;
  LAYER M1 ;
        RECT 63.085 31.415 63.335 34.945 ;
  LAYER M1 ;
        RECT 63.085 35.195 63.335 36.205 ;
  LAYER M1 ;
        RECT 63.085 37.295 63.335 40.825 ;
  LAYER M1 ;
        RECT 63.085 41.075 63.335 42.085 ;
  LAYER M1 ;
        RECT 63.085 43.175 63.335 46.705 ;
  LAYER M1 ;
        RECT 63.085 46.955 63.335 47.965 ;
  LAYER M1 ;
        RECT 63.085 49.055 63.335 52.585 ;
  LAYER M1 ;
        RECT 63.085 52.835 63.335 53.845 ;
  LAYER M1 ;
        RECT 63.085 54.935 63.335 55.945 ;
  LAYER M1 ;
        RECT 62.655 31.415 62.905 34.945 ;
  LAYER M1 ;
        RECT 62.655 37.295 62.905 40.825 ;
  LAYER M1 ;
        RECT 62.655 43.175 62.905 46.705 ;
  LAYER M1 ;
        RECT 62.655 49.055 62.905 52.585 ;
  LAYER M1 ;
        RECT 62.225 31.415 62.475 34.945 ;
  LAYER M1 ;
        RECT 62.225 35.195 62.475 36.205 ;
  LAYER M1 ;
        RECT 62.225 37.295 62.475 40.825 ;
  LAYER M1 ;
        RECT 62.225 41.075 62.475 42.085 ;
  LAYER M1 ;
        RECT 62.225 43.175 62.475 46.705 ;
  LAYER M1 ;
        RECT 62.225 46.955 62.475 47.965 ;
  LAYER M1 ;
        RECT 62.225 49.055 62.475 52.585 ;
  LAYER M1 ;
        RECT 62.225 52.835 62.475 53.845 ;
  LAYER M1 ;
        RECT 62.225 54.935 62.475 55.945 ;
  LAYER M1 ;
        RECT 61.795 31.415 62.045 34.945 ;
  LAYER M1 ;
        RECT 61.795 37.295 62.045 40.825 ;
  LAYER M1 ;
        RECT 61.795 43.175 62.045 46.705 ;
  LAYER M1 ;
        RECT 61.795 49.055 62.045 52.585 ;
  LAYER M1 ;
        RECT 61.365 31.415 61.615 34.945 ;
  LAYER M1 ;
        RECT 61.365 35.195 61.615 36.205 ;
  LAYER M1 ;
        RECT 61.365 37.295 61.615 40.825 ;
  LAYER M1 ;
        RECT 61.365 41.075 61.615 42.085 ;
  LAYER M1 ;
        RECT 61.365 43.175 61.615 46.705 ;
  LAYER M1 ;
        RECT 61.365 46.955 61.615 47.965 ;
  LAYER M1 ;
        RECT 61.365 49.055 61.615 52.585 ;
  LAYER M1 ;
        RECT 61.365 52.835 61.615 53.845 ;
  LAYER M1 ;
        RECT 61.365 54.935 61.615 55.945 ;
  LAYER M1 ;
        RECT 60.935 31.415 61.185 34.945 ;
  LAYER M1 ;
        RECT 60.935 37.295 61.185 40.825 ;
  LAYER M1 ;
        RECT 60.935 43.175 61.185 46.705 ;
  LAYER M1 ;
        RECT 60.935 49.055 61.185 52.585 ;
  LAYER M1 ;
        RECT 60.505 31.415 60.755 34.945 ;
  LAYER M1 ;
        RECT 60.505 35.195 60.755 36.205 ;
  LAYER M1 ;
        RECT 60.505 37.295 60.755 40.825 ;
  LAYER M1 ;
        RECT 60.505 41.075 60.755 42.085 ;
  LAYER M1 ;
        RECT 60.505 43.175 60.755 46.705 ;
  LAYER M1 ;
        RECT 60.505 46.955 60.755 47.965 ;
  LAYER M1 ;
        RECT 60.505 49.055 60.755 52.585 ;
  LAYER M1 ;
        RECT 60.505 52.835 60.755 53.845 ;
  LAYER M1 ;
        RECT 60.505 54.935 60.755 55.945 ;
  LAYER M1 ;
        RECT 60.075 31.415 60.325 34.945 ;
  LAYER M1 ;
        RECT 60.075 37.295 60.325 40.825 ;
  LAYER M1 ;
        RECT 60.075 43.175 60.325 46.705 ;
  LAYER M1 ;
        RECT 60.075 49.055 60.325 52.585 ;
  LAYER M1 ;
        RECT 59.645 31.415 59.895 34.945 ;
  LAYER M1 ;
        RECT 59.645 35.195 59.895 36.205 ;
  LAYER M1 ;
        RECT 59.645 37.295 59.895 40.825 ;
  LAYER M1 ;
        RECT 59.645 41.075 59.895 42.085 ;
  LAYER M1 ;
        RECT 59.645 43.175 59.895 46.705 ;
  LAYER M1 ;
        RECT 59.645 46.955 59.895 47.965 ;
  LAYER M1 ;
        RECT 59.645 49.055 59.895 52.585 ;
  LAYER M1 ;
        RECT 59.645 52.835 59.895 53.845 ;
  LAYER M1 ;
        RECT 59.645 54.935 59.895 55.945 ;
  LAYER M1 ;
        RECT 59.215 31.415 59.465 34.945 ;
  LAYER M1 ;
        RECT 59.215 37.295 59.465 40.825 ;
  LAYER M1 ;
        RECT 59.215 43.175 59.465 46.705 ;
  LAYER M1 ;
        RECT 59.215 49.055 59.465 52.585 ;
  LAYER M1 ;
        RECT 58.785 31.415 59.035 34.945 ;
  LAYER M1 ;
        RECT 58.785 35.195 59.035 36.205 ;
  LAYER M1 ;
        RECT 58.785 37.295 59.035 40.825 ;
  LAYER M1 ;
        RECT 58.785 41.075 59.035 42.085 ;
  LAYER M1 ;
        RECT 58.785 43.175 59.035 46.705 ;
  LAYER M1 ;
        RECT 58.785 46.955 59.035 47.965 ;
  LAYER M1 ;
        RECT 58.785 49.055 59.035 52.585 ;
  LAYER M1 ;
        RECT 58.785 52.835 59.035 53.845 ;
  LAYER M1 ;
        RECT 58.785 54.935 59.035 55.945 ;
  LAYER M1 ;
        RECT 58.355 31.415 58.605 34.945 ;
  LAYER M1 ;
        RECT 58.355 37.295 58.605 40.825 ;
  LAYER M1 ;
        RECT 58.355 43.175 58.605 46.705 ;
  LAYER M1 ;
        RECT 58.355 49.055 58.605 52.585 ;
  LAYER M1 ;
        RECT 57.925 31.415 58.175 34.945 ;
  LAYER M1 ;
        RECT 57.925 35.195 58.175 36.205 ;
  LAYER M1 ;
        RECT 57.925 37.295 58.175 40.825 ;
  LAYER M1 ;
        RECT 57.925 41.075 58.175 42.085 ;
  LAYER M1 ;
        RECT 57.925 43.175 58.175 46.705 ;
  LAYER M1 ;
        RECT 57.925 46.955 58.175 47.965 ;
  LAYER M1 ;
        RECT 57.925 49.055 58.175 52.585 ;
  LAYER M1 ;
        RECT 57.925 52.835 58.175 53.845 ;
  LAYER M1 ;
        RECT 57.925 54.935 58.175 55.945 ;
  LAYER M1 ;
        RECT 57.495 31.415 57.745 34.945 ;
  LAYER M1 ;
        RECT 57.495 37.295 57.745 40.825 ;
  LAYER M1 ;
        RECT 57.495 43.175 57.745 46.705 ;
  LAYER M1 ;
        RECT 57.495 49.055 57.745 52.585 ;
  LAYER M1 ;
        RECT 57.065 31.415 57.315 34.945 ;
  LAYER M1 ;
        RECT 57.065 35.195 57.315 36.205 ;
  LAYER M1 ;
        RECT 57.065 37.295 57.315 40.825 ;
  LAYER M1 ;
        RECT 57.065 41.075 57.315 42.085 ;
  LAYER M1 ;
        RECT 57.065 43.175 57.315 46.705 ;
  LAYER M1 ;
        RECT 57.065 46.955 57.315 47.965 ;
  LAYER M1 ;
        RECT 57.065 49.055 57.315 52.585 ;
  LAYER M1 ;
        RECT 57.065 52.835 57.315 53.845 ;
  LAYER M1 ;
        RECT 57.065 54.935 57.315 55.945 ;
  LAYER M1 ;
        RECT 56.635 31.415 56.885 34.945 ;
  LAYER M1 ;
        RECT 56.635 37.295 56.885 40.825 ;
  LAYER M1 ;
        RECT 56.635 43.175 56.885 46.705 ;
  LAYER M1 ;
        RECT 56.635 49.055 56.885 52.585 ;
  LAYER M1 ;
        RECT 56.205 31.415 56.455 34.945 ;
  LAYER M1 ;
        RECT 56.205 35.195 56.455 36.205 ;
  LAYER M1 ;
        RECT 56.205 37.295 56.455 40.825 ;
  LAYER M1 ;
        RECT 56.205 41.075 56.455 42.085 ;
  LAYER M1 ;
        RECT 56.205 43.175 56.455 46.705 ;
  LAYER M1 ;
        RECT 56.205 46.955 56.455 47.965 ;
  LAYER M1 ;
        RECT 56.205 49.055 56.455 52.585 ;
  LAYER M1 ;
        RECT 56.205 52.835 56.455 53.845 ;
  LAYER M1 ;
        RECT 56.205 54.935 56.455 55.945 ;
  LAYER M1 ;
        RECT 55.775 31.415 56.025 34.945 ;
  LAYER M1 ;
        RECT 55.775 37.295 56.025 40.825 ;
  LAYER M1 ;
        RECT 55.775 43.175 56.025 46.705 ;
  LAYER M1 ;
        RECT 55.775 49.055 56.025 52.585 ;
  LAYER M1 ;
        RECT 55.345 31.415 55.595 34.945 ;
  LAYER M1 ;
        RECT 55.345 35.195 55.595 36.205 ;
  LAYER M1 ;
        RECT 55.345 37.295 55.595 40.825 ;
  LAYER M1 ;
        RECT 55.345 41.075 55.595 42.085 ;
  LAYER M1 ;
        RECT 55.345 43.175 55.595 46.705 ;
  LAYER M1 ;
        RECT 55.345 46.955 55.595 47.965 ;
  LAYER M1 ;
        RECT 55.345 49.055 55.595 52.585 ;
  LAYER M1 ;
        RECT 55.345 52.835 55.595 53.845 ;
  LAYER M1 ;
        RECT 55.345 54.935 55.595 55.945 ;
  LAYER M1 ;
        RECT 54.915 31.415 55.165 34.945 ;
  LAYER M1 ;
        RECT 54.915 37.295 55.165 40.825 ;
  LAYER M1 ;
        RECT 54.915 43.175 55.165 46.705 ;
  LAYER M1 ;
        RECT 54.915 49.055 55.165 52.585 ;
  LAYER M1 ;
        RECT 54.485 31.415 54.735 34.945 ;
  LAYER M1 ;
        RECT 54.485 35.195 54.735 36.205 ;
  LAYER M1 ;
        RECT 54.485 37.295 54.735 40.825 ;
  LAYER M1 ;
        RECT 54.485 41.075 54.735 42.085 ;
  LAYER M1 ;
        RECT 54.485 43.175 54.735 46.705 ;
  LAYER M1 ;
        RECT 54.485 46.955 54.735 47.965 ;
  LAYER M1 ;
        RECT 54.485 49.055 54.735 52.585 ;
  LAYER M1 ;
        RECT 54.485 52.835 54.735 53.845 ;
  LAYER M1 ;
        RECT 54.485 54.935 54.735 55.945 ;
  LAYER M1 ;
        RECT 54.055 31.415 54.305 34.945 ;
  LAYER M1 ;
        RECT 54.055 37.295 54.305 40.825 ;
  LAYER M1 ;
        RECT 54.055 43.175 54.305 46.705 ;
  LAYER M1 ;
        RECT 54.055 49.055 54.305 52.585 ;
  LAYER M1 ;
        RECT 53.625 31.415 53.875 34.945 ;
  LAYER M1 ;
        RECT 53.625 35.195 53.875 36.205 ;
  LAYER M1 ;
        RECT 53.625 37.295 53.875 40.825 ;
  LAYER M1 ;
        RECT 53.625 41.075 53.875 42.085 ;
  LAYER M1 ;
        RECT 53.625 43.175 53.875 46.705 ;
  LAYER M1 ;
        RECT 53.625 46.955 53.875 47.965 ;
  LAYER M1 ;
        RECT 53.625 49.055 53.875 52.585 ;
  LAYER M1 ;
        RECT 53.625 52.835 53.875 53.845 ;
  LAYER M1 ;
        RECT 53.625 54.935 53.875 55.945 ;
  LAYER M1 ;
        RECT 53.195 31.415 53.445 34.945 ;
  LAYER M1 ;
        RECT 53.195 37.295 53.445 40.825 ;
  LAYER M1 ;
        RECT 53.195 43.175 53.445 46.705 ;
  LAYER M1 ;
        RECT 53.195 49.055 53.445 52.585 ;
  LAYER M1 ;
        RECT 52.765 31.415 53.015 34.945 ;
  LAYER M1 ;
        RECT 52.765 35.195 53.015 36.205 ;
  LAYER M1 ;
        RECT 52.765 37.295 53.015 40.825 ;
  LAYER M1 ;
        RECT 52.765 41.075 53.015 42.085 ;
  LAYER M1 ;
        RECT 52.765 43.175 53.015 46.705 ;
  LAYER M1 ;
        RECT 52.765 46.955 53.015 47.965 ;
  LAYER M1 ;
        RECT 52.765 49.055 53.015 52.585 ;
  LAYER M1 ;
        RECT 52.765 52.835 53.015 53.845 ;
  LAYER M1 ;
        RECT 52.765 54.935 53.015 55.945 ;
  LAYER M1 ;
        RECT 52.335 31.415 52.585 34.945 ;
  LAYER M1 ;
        RECT 52.335 37.295 52.585 40.825 ;
  LAYER M1 ;
        RECT 52.335 43.175 52.585 46.705 ;
  LAYER M1 ;
        RECT 52.335 49.055 52.585 52.585 ;
  LAYER M1 ;
        RECT 51.905 31.415 52.155 34.945 ;
  LAYER M1 ;
        RECT 51.905 35.195 52.155 36.205 ;
  LAYER M1 ;
        RECT 51.905 37.295 52.155 40.825 ;
  LAYER M1 ;
        RECT 51.905 41.075 52.155 42.085 ;
  LAYER M1 ;
        RECT 51.905 43.175 52.155 46.705 ;
  LAYER M1 ;
        RECT 51.905 46.955 52.155 47.965 ;
  LAYER M1 ;
        RECT 51.905 49.055 52.155 52.585 ;
  LAYER M1 ;
        RECT 51.905 52.835 52.155 53.845 ;
  LAYER M1 ;
        RECT 51.905 54.935 52.155 55.945 ;
  LAYER M1 ;
        RECT 51.475 31.415 51.725 34.945 ;
  LAYER M1 ;
        RECT 51.475 37.295 51.725 40.825 ;
  LAYER M1 ;
        RECT 51.475 43.175 51.725 46.705 ;
  LAYER M1 ;
        RECT 51.475 49.055 51.725 52.585 ;
  LAYER M1 ;
        RECT 51.045 31.415 51.295 34.945 ;
  LAYER M1 ;
        RECT 51.045 35.195 51.295 36.205 ;
  LAYER M1 ;
        RECT 51.045 37.295 51.295 40.825 ;
  LAYER M1 ;
        RECT 51.045 41.075 51.295 42.085 ;
  LAYER M1 ;
        RECT 51.045 43.175 51.295 46.705 ;
  LAYER M1 ;
        RECT 51.045 46.955 51.295 47.965 ;
  LAYER M1 ;
        RECT 51.045 49.055 51.295 52.585 ;
  LAYER M1 ;
        RECT 51.045 52.835 51.295 53.845 ;
  LAYER M1 ;
        RECT 51.045 54.935 51.295 55.945 ;
  LAYER M1 ;
        RECT 50.615 31.415 50.865 34.945 ;
  LAYER M1 ;
        RECT 50.615 37.295 50.865 40.825 ;
  LAYER M1 ;
        RECT 50.615 43.175 50.865 46.705 ;
  LAYER M1 ;
        RECT 50.615 49.055 50.865 52.585 ;
  LAYER M1 ;
        RECT 50.185 31.415 50.435 34.945 ;
  LAYER M1 ;
        RECT 50.185 35.195 50.435 36.205 ;
  LAYER M1 ;
        RECT 50.185 37.295 50.435 40.825 ;
  LAYER M1 ;
        RECT 50.185 41.075 50.435 42.085 ;
  LAYER M1 ;
        RECT 50.185 43.175 50.435 46.705 ;
  LAYER M1 ;
        RECT 50.185 46.955 50.435 47.965 ;
  LAYER M1 ;
        RECT 50.185 49.055 50.435 52.585 ;
  LAYER M1 ;
        RECT 50.185 52.835 50.435 53.845 ;
  LAYER M1 ;
        RECT 50.185 54.935 50.435 55.945 ;
  LAYER M1 ;
        RECT 49.755 31.415 50.005 34.945 ;
  LAYER M1 ;
        RECT 49.755 37.295 50.005 40.825 ;
  LAYER M1 ;
        RECT 49.755 43.175 50.005 46.705 ;
  LAYER M1 ;
        RECT 49.755 49.055 50.005 52.585 ;
  LAYER M1 ;
        RECT 49.325 31.415 49.575 34.945 ;
  LAYER M1 ;
        RECT 49.325 35.195 49.575 36.205 ;
  LAYER M1 ;
        RECT 49.325 37.295 49.575 40.825 ;
  LAYER M1 ;
        RECT 49.325 41.075 49.575 42.085 ;
  LAYER M1 ;
        RECT 49.325 43.175 49.575 46.705 ;
  LAYER M1 ;
        RECT 49.325 46.955 49.575 47.965 ;
  LAYER M1 ;
        RECT 49.325 49.055 49.575 52.585 ;
  LAYER M1 ;
        RECT 49.325 52.835 49.575 53.845 ;
  LAYER M1 ;
        RECT 49.325 54.935 49.575 55.945 ;
  LAYER M1 ;
        RECT 48.895 31.415 49.145 34.945 ;
  LAYER M1 ;
        RECT 48.895 37.295 49.145 40.825 ;
  LAYER M1 ;
        RECT 48.895 43.175 49.145 46.705 ;
  LAYER M1 ;
        RECT 48.895 49.055 49.145 52.585 ;
  LAYER M1 ;
        RECT 48.465 31.415 48.715 34.945 ;
  LAYER M1 ;
        RECT 48.465 35.195 48.715 36.205 ;
  LAYER M1 ;
        RECT 48.465 37.295 48.715 40.825 ;
  LAYER M1 ;
        RECT 48.465 41.075 48.715 42.085 ;
  LAYER M1 ;
        RECT 48.465 43.175 48.715 46.705 ;
  LAYER M1 ;
        RECT 48.465 46.955 48.715 47.965 ;
  LAYER M1 ;
        RECT 48.465 49.055 48.715 52.585 ;
  LAYER M1 ;
        RECT 48.465 52.835 48.715 53.845 ;
  LAYER M1 ;
        RECT 48.465 54.935 48.715 55.945 ;
  LAYER M1 ;
        RECT 48.035 31.415 48.285 34.945 ;
  LAYER M1 ;
        RECT 48.035 37.295 48.285 40.825 ;
  LAYER M1 ;
        RECT 48.035 43.175 48.285 46.705 ;
  LAYER M1 ;
        RECT 48.035 49.055 48.285 52.585 ;
  LAYER M1 ;
        RECT 47.605 31.415 47.855 34.945 ;
  LAYER M1 ;
        RECT 47.605 35.195 47.855 36.205 ;
  LAYER M1 ;
        RECT 47.605 37.295 47.855 40.825 ;
  LAYER M1 ;
        RECT 47.605 41.075 47.855 42.085 ;
  LAYER M1 ;
        RECT 47.605 43.175 47.855 46.705 ;
  LAYER M1 ;
        RECT 47.605 46.955 47.855 47.965 ;
  LAYER M1 ;
        RECT 47.605 49.055 47.855 52.585 ;
  LAYER M1 ;
        RECT 47.605 52.835 47.855 53.845 ;
  LAYER M1 ;
        RECT 47.605 54.935 47.855 55.945 ;
  LAYER M1 ;
        RECT 47.175 31.415 47.425 34.945 ;
  LAYER M1 ;
        RECT 47.175 37.295 47.425 40.825 ;
  LAYER M1 ;
        RECT 47.175 43.175 47.425 46.705 ;
  LAYER M1 ;
        RECT 47.175 49.055 47.425 52.585 ;
  LAYER M1 ;
        RECT 46.745 31.415 46.995 34.945 ;
  LAYER M1 ;
        RECT 46.745 35.195 46.995 36.205 ;
  LAYER M1 ;
        RECT 46.745 37.295 46.995 40.825 ;
  LAYER M1 ;
        RECT 46.745 41.075 46.995 42.085 ;
  LAYER M1 ;
        RECT 46.745 43.175 46.995 46.705 ;
  LAYER M1 ;
        RECT 46.745 46.955 46.995 47.965 ;
  LAYER M1 ;
        RECT 46.745 49.055 46.995 52.585 ;
  LAYER M1 ;
        RECT 46.745 52.835 46.995 53.845 ;
  LAYER M1 ;
        RECT 46.745 54.935 46.995 55.945 ;
  LAYER M1 ;
        RECT 46.315 31.415 46.565 34.945 ;
  LAYER M1 ;
        RECT 46.315 37.295 46.565 40.825 ;
  LAYER M1 ;
        RECT 46.315 43.175 46.565 46.705 ;
  LAYER M1 ;
        RECT 46.315 49.055 46.565 52.585 ;
  LAYER M1 ;
        RECT 45.885 31.415 46.135 34.945 ;
  LAYER M1 ;
        RECT 45.885 35.195 46.135 36.205 ;
  LAYER M1 ;
        RECT 45.885 37.295 46.135 40.825 ;
  LAYER M1 ;
        RECT 45.885 41.075 46.135 42.085 ;
  LAYER M1 ;
        RECT 45.885 43.175 46.135 46.705 ;
  LAYER M1 ;
        RECT 45.885 46.955 46.135 47.965 ;
  LAYER M1 ;
        RECT 45.885 49.055 46.135 52.585 ;
  LAYER M1 ;
        RECT 45.885 52.835 46.135 53.845 ;
  LAYER M1 ;
        RECT 45.885 54.935 46.135 55.945 ;
  LAYER M1 ;
        RECT 45.455 31.415 45.705 34.945 ;
  LAYER M1 ;
        RECT 45.455 37.295 45.705 40.825 ;
  LAYER M1 ;
        RECT 45.455 43.175 45.705 46.705 ;
  LAYER M1 ;
        RECT 45.455 49.055 45.705 52.585 ;
  LAYER M1 ;
        RECT 45.025 31.415 45.275 34.945 ;
  LAYER M1 ;
        RECT 45.025 35.195 45.275 36.205 ;
  LAYER M1 ;
        RECT 45.025 37.295 45.275 40.825 ;
  LAYER M1 ;
        RECT 45.025 41.075 45.275 42.085 ;
  LAYER M1 ;
        RECT 45.025 43.175 45.275 46.705 ;
  LAYER M1 ;
        RECT 45.025 46.955 45.275 47.965 ;
  LAYER M1 ;
        RECT 45.025 49.055 45.275 52.585 ;
  LAYER M1 ;
        RECT 45.025 52.835 45.275 53.845 ;
  LAYER M1 ;
        RECT 45.025 54.935 45.275 55.945 ;
  LAYER M1 ;
        RECT 44.595 31.415 44.845 34.945 ;
  LAYER M1 ;
        RECT 44.595 37.295 44.845 40.825 ;
  LAYER M1 ;
        RECT 44.595 43.175 44.845 46.705 ;
  LAYER M1 ;
        RECT 44.595 49.055 44.845 52.585 ;
  LAYER M1 ;
        RECT 44.165 31.415 44.415 34.945 ;
  LAYER M1 ;
        RECT 44.165 35.195 44.415 36.205 ;
  LAYER M1 ;
        RECT 44.165 37.295 44.415 40.825 ;
  LAYER M1 ;
        RECT 44.165 41.075 44.415 42.085 ;
  LAYER M1 ;
        RECT 44.165 43.175 44.415 46.705 ;
  LAYER M1 ;
        RECT 44.165 46.955 44.415 47.965 ;
  LAYER M1 ;
        RECT 44.165 49.055 44.415 52.585 ;
  LAYER M1 ;
        RECT 44.165 52.835 44.415 53.845 ;
  LAYER M1 ;
        RECT 44.165 54.935 44.415 55.945 ;
  LAYER M1 ;
        RECT 43.735 31.415 43.985 34.945 ;
  LAYER M1 ;
        RECT 43.735 37.295 43.985 40.825 ;
  LAYER M1 ;
        RECT 43.735 43.175 43.985 46.705 ;
  LAYER M1 ;
        RECT 43.735 49.055 43.985 52.585 ;
  LAYER M1 ;
        RECT 43.305 31.415 43.555 34.945 ;
  LAYER M1 ;
        RECT 43.305 35.195 43.555 36.205 ;
  LAYER M1 ;
        RECT 43.305 37.295 43.555 40.825 ;
  LAYER M1 ;
        RECT 43.305 41.075 43.555 42.085 ;
  LAYER M1 ;
        RECT 43.305 43.175 43.555 46.705 ;
  LAYER M1 ;
        RECT 43.305 46.955 43.555 47.965 ;
  LAYER M1 ;
        RECT 43.305 49.055 43.555 52.585 ;
  LAYER M1 ;
        RECT 43.305 52.835 43.555 53.845 ;
  LAYER M1 ;
        RECT 43.305 54.935 43.555 55.945 ;
  LAYER M1 ;
        RECT 42.875 31.415 43.125 34.945 ;
  LAYER M1 ;
        RECT 42.875 37.295 43.125 40.825 ;
  LAYER M1 ;
        RECT 42.875 43.175 43.125 46.705 ;
  LAYER M1 ;
        RECT 42.875 49.055 43.125 52.585 ;
  LAYER M1 ;
        RECT 42.445 31.415 42.695 34.945 ;
  LAYER M1 ;
        RECT 42.445 35.195 42.695 36.205 ;
  LAYER M1 ;
        RECT 42.445 37.295 42.695 40.825 ;
  LAYER M1 ;
        RECT 42.445 41.075 42.695 42.085 ;
  LAYER M1 ;
        RECT 42.445 43.175 42.695 46.705 ;
  LAYER M1 ;
        RECT 42.445 46.955 42.695 47.965 ;
  LAYER M1 ;
        RECT 42.445 49.055 42.695 52.585 ;
  LAYER M1 ;
        RECT 42.445 52.835 42.695 53.845 ;
  LAYER M1 ;
        RECT 42.445 54.935 42.695 55.945 ;
  LAYER M1 ;
        RECT 42.015 31.415 42.265 34.945 ;
  LAYER M1 ;
        RECT 42.015 37.295 42.265 40.825 ;
  LAYER M1 ;
        RECT 42.015 43.175 42.265 46.705 ;
  LAYER M1 ;
        RECT 42.015 49.055 42.265 52.585 ;
  LAYER M1 ;
        RECT 41.585 31.415 41.835 34.945 ;
  LAYER M1 ;
        RECT 41.585 35.195 41.835 36.205 ;
  LAYER M1 ;
        RECT 41.585 37.295 41.835 40.825 ;
  LAYER M1 ;
        RECT 41.585 41.075 41.835 42.085 ;
  LAYER M1 ;
        RECT 41.585 43.175 41.835 46.705 ;
  LAYER M1 ;
        RECT 41.585 46.955 41.835 47.965 ;
  LAYER M1 ;
        RECT 41.585 49.055 41.835 52.585 ;
  LAYER M1 ;
        RECT 41.585 52.835 41.835 53.845 ;
  LAYER M1 ;
        RECT 41.585 54.935 41.835 55.945 ;
  LAYER M1 ;
        RECT 41.155 31.415 41.405 34.945 ;
  LAYER M1 ;
        RECT 41.155 37.295 41.405 40.825 ;
  LAYER M1 ;
        RECT 41.155 43.175 41.405 46.705 ;
  LAYER M1 ;
        RECT 41.155 49.055 41.405 52.585 ;
  LAYER M1 ;
        RECT 40.725 31.415 40.975 34.945 ;
  LAYER M1 ;
        RECT 40.725 35.195 40.975 36.205 ;
  LAYER M1 ;
        RECT 40.725 37.295 40.975 40.825 ;
  LAYER M1 ;
        RECT 40.725 41.075 40.975 42.085 ;
  LAYER M1 ;
        RECT 40.725 43.175 40.975 46.705 ;
  LAYER M1 ;
        RECT 40.725 46.955 40.975 47.965 ;
  LAYER M1 ;
        RECT 40.725 49.055 40.975 52.585 ;
  LAYER M1 ;
        RECT 40.725 52.835 40.975 53.845 ;
  LAYER M1 ;
        RECT 40.725 54.935 40.975 55.945 ;
  LAYER M1 ;
        RECT 40.295 31.415 40.545 34.945 ;
  LAYER M1 ;
        RECT 40.295 37.295 40.545 40.825 ;
  LAYER M1 ;
        RECT 40.295 43.175 40.545 46.705 ;
  LAYER M1 ;
        RECT 40.295 49.055 40.545 52.585 ;
  LAYER M1 ;
        RECT 39.865 31.415 40.115 34.945 ;
  LAYER M1 ;
        RECT 39.865 35.195 40.115 36.205 ;
  LAYER M1 ;
        RECT 39.865 37.295 40.115 40.825 ;
  LAYER M1 ;
        RECT 39.865 41.075 40.115 42.085 ;
  LAYER M1 ;
        RECT 39.865 43.175 40.115 46.705 ;
  LAYER M1 ;
        RECT 39.865 46.955 40.115 47.965 ;
  LAYER M1 ;
        RECT 39.865 49.055 40.115 52.585 ;
  LAYER M1 ;
        RECT 39.865 52.835 40.115 53.845 ;
  LAYER M1 ;
        RECT 39.865 54.935 40.115 55.945 ;
  LAYER M1 ;
        RECT 39.435 31.415 39.685 34.945 ;
  LAYER M1 ;
        RECT 39.435 37.295 39.685 40.825 ;
  LAYER M1 ;
        RECT 39.435 43.175 39.685 46.705 ;
  LAYER M1 ;
        RECT 39.435 49.055 39.685 52.585 ;
  LAYER M1 ;
        RECT 39.005 31.415 39.255 34.945 ;
  LAYER M1 ;
        RECT 39.005 35.195 39.255 36.205 ;
  LAYER M1 ;
        RECT 39.005 37.295 39.255 40.825 ;
  LAYER M1 ;
        RECT 39.005 41.075 39.255 42.085 ;
  LAYER M1 ;
        RECT 39.005 43.175 39.255 46.705 ;
  LAYER M1 ;
        RECT 39.005 46.955 39.255 47.965 ;
  LAYER M1 ;
        RECT 39.005 49.055 39.255 52.585 ;
  LAYER M1 ;
        RECT 39.005 52.835 39.255 53.845 ;
  LAYER M1 ;
        RECT 39.005 54.935 39.255 55.945 ;
  LAYER M1 ;
        RECT 38.575 31.415 38.825 34.945 ;
  LAYER M1 ;
        RECT 38.575 37.295 38.825 40.825 ;
  LAYER M1 ;
        RECT 38.575 43.175 38.825 46.705 ;
  LAYER M1 ;
        RECT 38.575 49.055 38.825 52.585 ;
  LAYER M1 ;
        RECT 38.145 31.415 38.395 34.945 ;
  LAYER M1 ;
        RECT 38.145 35.195 38.395 36.205 ;
  LAYER M1 ;
        RECT 38.145 37.295 38.395 40.825 ;
  LAYER M1 ;
        RECT 38.145 41.075 38.395 42.085 ;
  LAYER M1 ;
        RECT 38.145 43.175 38.395 46.705 ;
  LAYER M1 ;
        RECT 38.145 46.955 38.395 47.965 ;
  LAYER M1 ;
        RECT 38.145 49.055 38.395 52.585 ;
  LAYER M1 ;
        RECT 38.145 52.835 38.395 53.845 ;
  LAYER M1 ;
        RECT 38.145 54.935 38.395 55.945 ;
  LAYER M1 ;
        RECT 37.715 31.415 37.965 34.945 ;
  LAYER M1 ;
        RECT 37.715 37.295 37.965 40.825 ;
  LAYER M1 ;
        RECT 37.715 43.175 37.965 46.705 ;
  LAYER M1 ;
        RECT 37.715 49.055 37.965 52.585 ;
  LAYER M1 ;
        RECT 37.285 31.415 37.535 34.945 ;
  LAYER M1 ;
        RECT 37.285 35.195 37.535 36.205 ;
  LAYER M1 ;
        RECT 37.285 37.295 37.535 40.825 ;
  LAYER M1 ;
        RECT 37.285 41.075 37.535 42.085 ;
  LAYER M1 ;
        RECT 37.285 43.175 37.535 46.705 ;
  LAYER M1 ;
        RECT 37.285 46.955 37.535 47.965 ;
  LAYER M1 ;
        RECT 37.285 49.055 37.535 52.585 ;
  LAYER M1 ;
        RECT 37.285 52.835 37.535 53.845 ;
  LAYER M1 ;
        RECT 37.285 54.935 37.535 55.945 ;
  LAYER M1 ;
        RECT 36.855 31.415 37.105 34.945 ;
  LAYER M1 ;
        RECT 36.855 37.295 37.105 40.825 ;
  LAYER M1 ;
        RECT 36.855 43.175 37.105 46.705 ;
  LAYER M1 ;
        RECT 36.855 49.055 37.105 52.585 ;
  LAYER M1 ;
        RECT 36.425 31.415 36.675 34.945 ;
  LAYER M1 ;
        RECT 36.425 35.195 36.675 36.205 ;
  LAYER M1 ;
        RECT 36.425 37.295 36.675 40.825 ;
  LAYER M1 ;
        RECT 36.425 41.075 36.675 42.085 ;
  LAYER M1 ;
        RECT 36.425 43.175 36.675 46.705 ;
  LAYER M1 ;
        RECT 36.425 46.955 36.675 47.965 ;
  LAYER M1 ;
        RECT 36.425 49.055 36.675 52.585 ;
  LAYER M1 ;
        RECT 36.425 52.835 36.675 53.845 ;
  LAYER M1 ;
        RECT 36.425 54.935 36.675 55.945 ;
  LAYER M1 ;
        RECT 35.995 31.415 36.245 34.945 ;
  LAYER M1 ;
        RECT 35.995 37.295 36.245 40.825 ;
  LAYER M1 ;
        RECT 35.995 43.175 36.245 46.705 ;
  LAYER M1 ;
        RECT 35.995 49.055 36.245 52.585 ;
  LAYER M1 ;
        RECT 35.565 31.415 35.815 34.945 ;
  LAYER M1 ;
        RECT 35.565 35.195 35.815 36.205 ;
  LAYER M1 ;
        RECT 35.565 37.295 35.815 40.825 ;
  LAYER M1 ;
        RECT 35.565 41.075 35.815 42.085 ;
  LAYER M1 ;
        RECT 35.565 43.175 35.815 46.705 ;
  LAYER M1 ;
        RECT 35.565 46.955 35.815 47.965 ;
  LAYER M1 ;
        RECT 35.565 49.055 35.815 52.585 ;
  LAYER M1 ;
        RECT 35.565 52.835 35.815 53.845 ;
  LAYER M1 ;
        RECT 35.565 54.935 35.815 55.945 ;
  LAYER M1 ;
        RECT 35.135 31.415 35.385 34.945 ;
  LAYER M1 ;
        RECT 35.135 37.295 35.385 40.825 ;
  LAYER M1 ;
        RECT 35.135 43.175 35.385 46.705 ;
  LAYER M1 ;
        RECT 35.135 49.055 35.385 52.585 ;
  LAYER M1 ;
        RECT 34.705 31.415 34.955 34.945 ;
  LAYER M1 ;
        RECT 34.705 35.195 34.955 36.205 ;
  LAYER M1 ;
        RECT 34.705 37.295 34.955 40.825 ;
  LAYER M1 ;
        RECT 34.705 41.075 34.955 42.085 ;
  LAYER M1 ;
        RECT 34.705 43.175 34.955 46.705 ;
  LAYER M1 ;
        RECT 34.705 46.955 34.955 47.965 ;
  LAYER M1 ;
        RECT 34.705 49.055 34.955 52.585 ;
  LAYER M1 ;
        RECT 34.705 52.835 34.955 53.845 ;
  LAYER M1 ;
        RECT 34.705 54.935 34.955 55.945 ;
  LAYER M1 ;
        RECT 34.275 31.415 34.525 34.945 ;
  LAYER M1 ;
        RECT 34.275 37.295 34.525 40.825 ;
  LAYER M1 ;
        RECT 34.275 43.175 34.525 46.705 ;
  LAYER M1 ;
        RECT 34.275 49.055 34.525 52.585 ;
  LAYER M2 ;
        RECT 34.66 31.36 65.96 31.64 ;
  LAYER M2 ;
        RECT 34.66 35.56 65.96 35.84 ;
  LAYER M2 ;
        RECT 34.23 31.78 66.39 32.06 ;
  LAYER M2 ;
        RECT 34.66 37.24 65.96 37.52 ;
  LAYER M2 ;
        RECT 34.66 41.44 65.96 41.72 ;
  LAYER M2 ;
        RECT 34.23 37.66 66.39 37.94 ;
  LAYER M2 ;
        RECT 34.66 43.12 65.96 43.4 ;
  LAYER M2 ;
        RECT 34.66 47.32 65.96 47.6 ;
  LAYER M2 ;
        RECT 34.23 43.54 66.39 43.82 ;
  LAYER M2 ;
        RECT 34.66 49 65.96 49.28 ;
  LAYER M2 ;
        RECT 34.66 53.2 65.96 53.48 ;
  LAYER M2 ;
        RECT 34.66 55.3 65.96 55.58 ;
  LAYER M2 ;
        RECT 34.23 49.42 66.39 49.7 ;
  LAYER M3 ;
        RECT 50.6 31.34 50.88 49.3 ;
  LAYER M3 ;
        RECT 50.17 35.54 50.45 53.5 ;
  LAYER M3 ;
        RECT 49.74 31.76 50.02 55.6 ;
  LAYER M1 ;
        RECT 34.705 0.335 34.955 3.865 ;
  LAYER M1 ;
        RECT 34.705 4.115 34.955 5.125 ;
  LAYER M1 ;
        RECT 34.705 6.215 34.955 9.745 ;
  LAYER M1 ;
        RECT 34.705 9.995 34.955 11.005 ;
  LAYER M1 ;
        RECT 34.705 12.095 34.955 15.625 ;
  LAYER M1 ;
        RECT 34.705 15.875 34.955 16.885 ;
  LAYER M1 ;
        RECT 34.705 17.975 34.955 21.505 ;
  LAYER M1 ;
        RECT 34.705 21.755 34.955 22.765 ;
  LAYER M1 ;
        RECT 34.705 23.855 34.955 27.385 ;
  LAYER M1 ;
        RECT 34.705 27.635 34.955 28.645 ;
  LAYER M1 ;
        RECT 34.705 29.735 34.955 30.745 ;
  LAYER M1 ;
        RECT 34.275 0.335 34.525 3.865 ;
  LAYER M1 ;
        RECT 34.275 6.215 34.525 9.745 ;
  LAYER M1 ;
        RECT 34.275 12.095 34.525 15.625 ;
  LAYER M1 ;
        RECT 34.275 17.975 34.525 21.505 ;
  LAYER M1 ;
        RECT 34.275 23.855 34.525 27.385 ;
  LAYER M1 ;
        RECT 35.135 0.335 35.385 3.865 ;
  LAYER M1 ;
        RECT 35.135 6.215 35.385 9.745 ;
  LAYER M1 ;
        RECT 35.135 12.095 35.385 15.625 ;
  LAYER M1 ;
        RECT 35.135 17.975 35.385 21.505 ;
  LAYER M1 ;
        RECT 35.135 23.855 35.385 27.385 ;
  LAYER M1 ;
        RECT 35.565 0.335 35.815 3.865 ;
  LAYER M1 ;
        RECT 35.565 4.115 35.815 5.125 ;
  LAYER M1 ;
        RECT 35.565 6.215 35.815 9.745 ;
  LAYER M1 ;
        RECT 35.565 9.995 35.815 11.005 ;
  LAYER M1 ;
        RECT 35.565 12.095 35.815 15.625 ;
  LAYER M1 ;
        RECT 35.565 15.875 35.815 16.885 ;
  LAYER M1 ;
        RECT 35.565 17.975 35.815 21.505 ;
  LAYER M1 ;
        RECT 35.565 21.755 35.815 22.765 ;
  LAYER M1 ;
        RECT 35.565 23.855 35.815 27.385 ;
  LAYER M1 ;
        RECT 35.565 27.635 35.815 28.645 ;
  LAYER M1 ;
        RECT 35.565 29.735 35.815 30.745 ;
  LAYER M1 ;
        RECT 35.995 0.335 36.245 3.865 ;
  LAYER M1 ;
        RECT 35.995 6.215 36.245 9.745 ;
  LAYER M1 ;
        RECT 35.995 12.095 36.245 15.625 ;
  LAYER M1 ;
        RECT 35.995 17.975 36.245 21.505 ;
  LAYER M1 ;
        RECT 35.995 23.855 36.245 27.385 ;
  LAYER M1 ;
        RECT 36.425 0.335 36.675 3.865 ;
  LAYER M1 ;
        RECT 36.425 4.115 36.675 5.125 ;
  LAYER M1 ;
        RECT 36.425 6.215 36.675 9.745 ;
  LAYER M1 ;
        RECT 36.425 9.995 36.675 11.005 ;
  LAYER M1 ;
        RECT 36.425 12.095 36.675 15.625 ;
  LAYER M1 ;
        RECT 36.425 15.875 36.675 16.885 ;
  LAYER M1 ;
        RECT 36.425 17.975 36.675 21.505 ;
  LAYER M1 ;
        RECT 36.425 21.755 36.675 22.765 ;
  LAYER M1 ;
        RECT 36.425 23.855 36.675 27.385 ;
  LAYER M1 ;
        RECT 36.425 27.635 36.675 28.645 ;
  LAYER M1 ;
        RECT 36.425 29.735 36.675 30.745 ;
  LAYER M1 ;
        RECT 36.855 0.335 37.105 3.865 ;
  LAYER M1 ;
        RECT 36.855 6.215 37.105 9.745 ;
  LAYER M1 ;
        RECT 36.855 12.095 37.105 15.625 ;
  LAYER M1 ;
        RECT 36.855 17.975 37.105 21.505 ;
  LAYER M1 ;
        RECT 36.855 23.855 37.105 27.385 ;
  LAYER M1 ;
        RECT 37.285 0.335 37.535 3.865 ;
  LAYER M1 ;
        RECT 37.285 4.115 37.535 5.125 ;
  LAYER M1 ;
        RECT 37.285 6.215 37.535 9.745 ;
  LAYER M1 ;
        RECT 37.285 9.995 37.535 11.005 ;
  LAYER M1 ;
        RECT 37.285 12.095 37.535 15.625 ;
  LAYER M1 ;
        RECT 37.285 15.875 37.535 16.885 ;
  LAYER M1 ;
        RECT 37.285 17.975 37.535 21.505 ;
  LAYER M1 ;
        RECT 37.285 21.755 37.535 22.765 ;
  LAYER M1 ;
        RECT 37.285 23.855 37.535 27.385 ;
  LAYER M1 ;
        RECT 37.285 27.635 37.535 28.645 ;
  LAYER M1 ;
        RECT 37.285 29.735 37.535 30.745 ;
  LAYER M1 ;
        RECT 37.715 0.335 37.965 3.865 ;
  LAYER M1 ;
        RECT 37.715 6.215 37.965 9.745 ;
  LAYER M1 ;
        RECT 37.715 12.095 37.965 15.625 ;
  LAYER M1 ;
        RECT 37.715 17.975 37.965 21.505 ;
  LAYER M1 ;
        RECT 37.715 23.855 37.965 27.385 ;
  LAYER M1 ;
        RECT 38.145 0.335 38.395 3.865 ;
  LAYER M1 ;
        RECT 38.145 4.115 38.395 5.125 ;
  LAYER M1 ;
        RECT 38.145 6.215 38.395 9.745 ;
  LAYER M1 ;
        RECT 38.145 9.995 38.395 11.005 ;
  LAYER M1 ;
        RECT 38.145 12.095 38.395 15.625 ;
  LAYER M1 ;
        RECT 38.145 15.875 38.395 16.885 ;
  LAYER M1 ;
        RECT 38.145 17.975 38.395 21.505 ;
  LAYER M1 ;
        RECT 38.145 21.755 38.395 22.765 ;
  LAYER M1 ;
        RECT 38.145 23.855 38.395 27.385 ;
  LAYER M1 ;
        RECT 38.145 27.635 38.395 28.645 ;
  LAYER M1 ;
        RECT 38.145 29.735 38.395 30.745 ;
  LAYER M1 ;
        RECT 38.575 0.335 38.825 3.865 ;
  LAYER M1 ;
        RECT 38.575 6.215 38.825 9.745 ;
  LAYER M1 ;
        RECT 38.575 12.095 38.825 15.625 ;
  LAYER M1 ;
        RECT 38.575 17.975 38.825 21.505 ;
  LAYER M1 ;
        RECT 38.575 23.855 38.825 27.385 ;
  LAYER M1 ;
        RECT 39.005 0.335 39.255 3.865 ;
  LAYER M1 ;
        RECT 39.005 4.115 39.255 5.125 ;
  LAYER M1 ;
        RECT 39.005 6.215 39.255 9.745 ;
  LAYER M1 ;
        RECT 39.005 9.995 39.255 11.005 ;
  LAYER M1 ;
        RECT 39.005 12.095 39.255 15.625 ;
  LAYER M1 ;
        RECT 39.005 15.875 39.255 16.885 ;
  LAYER M1 ;
        RECT 39.005 17.975 39.255 21.505 ;
  LAYER M1 ;
        RECT 39.005 21.755 39.255 22.765 ;
  LAYER M1 ;
        RECT 39.005 23.855 39.255 27.385 ;
  LAYER M1 ;
        RECT 39.005 27.635 39.255 28.645 ;
  LAYER M1 ;
        RECT 39.005 29.735 39.255 30.745 ;
  LAYER M1 ;
        RECT 39.435 0.335 39.685 3.865 ;
  LAYER M1 ;
        RECT 39.435 6.215 39.685 9.745 ;
  LAYER M1 ;
        RECT 39.435 12.095 39.685 15.625 ;
  LAYER M1 ;
        RECT 39.435 17.975 39.685 21.505 ;
  LAYER M1 ;
        RECT 39.435 23.855 39.685 27.385 ;
  LAYER M1 ;
        RECT 39.865 0.335 40.115 3.865 ;
  LAYER M1 ;
        RECT 39.865 4.115 40.115 5.125 ;
  LAYER M1 ;
        RECT 39.865 6.215 40.115 9.745 ;
  LAYER M1 ;
        RECT 39.865 9.995 40.115 11.005 ;
  LAYER M1 ;
        RECT 39.865 12.095 40.115 15.625 ;
  LAYER M1 ;
        RECT 39.865 15.875 40.115 16.885 ;
  LAYER M1 ;
        RECT 39.865 17.975 40.115 21.505 ;
  LAYER M1 ;
        RECT 39.865 21.755 40.115 22.765 ;
  LAYER M1 ;
        RECT 39.865 23.855 40.115 27.385 ;
  LAYER M1 ;
        RECT 39.865 27.635 40.115 28.645 ;
  LAYER M1 ;
        RECT 39.865 29.735 40.115 30.745 ;
  LAYER M1 ;
        RECT 40.295 0.335 40.545 3.865 ;
  LAYER M1 ;
        RECT 40.295 6.215 40.545 9.745 ;
  LAYER M1 ;
        RECT 40.295 12.095 40.545 15.625 ;
  LAYER M1 ;
        RECT 40.295 17.975 40.545 21.505 ;
  LAYER M1 ;
        RECT 40.295 23.855 40.545 27.385 ;
  LAYER M1 ;
        RECT 40.725 0.335 40.975 3.865 ;
  LAYER M1 ;
        RECT 40.725 4.115 40.975 5.125 ;
  LAYER M1 ;
        RECT 40.725 6.215 40.975 9.745 ;
  LAYER M1 ;
        RECT 40.725 9.995 40.975 11.005 ;
  LAYER M1 ;
        RECT 40.725 12.095 40.975 15.625 ;
  LAYER M1 ;
        RECT 40.725 15.875 40.975 16.885 ;
  LAYER M1 ;
        RECT 40.725 17.975 40.975 21.505 ;
  LAYER M1 ;
        RECT 40.725 21.755 40.975 22.765 ;
  LAYER M1 ;
        RECT 40.725 23.855 40.975 27.385 ;
  LAYER M1 ;
        RECT 40.725 27.635 40.975 28.645 ;
  LAYER M1 ;
        RECT 40.725 29.735 40.975 30.745 ;
  LAYER M1 ;
        RECT 41.155 0.335 41.405 3.865 ;
  LAYER M1 ;
        RECT 41.155 6.215 41.405 9.745 ;
  LAYER M1 ;
        RECT 41.155 12.095 41.405 15.625 ;
  LAYER M1 ;
        RECT 41.155 17.975 41.405 21.505 ;
  LAYER M1 ;
        RECT 41.155 23.855 41.405 27.385 ;
  LAYER M1 ;
        RECT 41.585 0.335 41.835 3.865 ;
  LAYER M1 ;
        RECT 41.585 4.115 41.835 5.125 ;
  LAYER M1 ;
        RECT 41.585 6.215 41.835 9.745 ;
  LAYER M1 ;
        RECT 41.585 9.995 41.835 11.005 ;
  LAYER M1 ;
        RECT 41.585 12.095 41.835 15.625 ;
  LAYER M1 ;
        RECT 41.585 15.875 41.835 16.885 ;
  LAYER M1 ;
        RECT 41.585 17.975 41.835 21.505 ;
  LAYER M1 ;
        RECT 41.585 21.755 41.835 22.765 ;
  LAYER M1 ;
        RECT 41.585 23.855 41.835 27.385 ;
  LAYER M1 ;
        RECT 41.585 27.635 41.835 28.645 ;
  LAYER M1 ;
        RECT 41.585 29.735 41.835 30.745 ;
  LAYER M1 ;
        RECT 42.015 0.335 42.265 3.865 ;
  LAYER M1 ;
        RECT 42.015 6.215 42.265 9.745 ;
  LAYER M1 ;
        RECT 42.015 12.095 42.265 15.625 ;
  LAYER M1 ;
        RECT 42.015 17.975 42.265 21.505 ;
  LAYER M1 ;
        RECT 42.015 23.855 42.265 27.385 ;
  LAYER M1 ;
        RECT 42.445 0.335 42.695 3.865 ;
  LAYER M1 ;
        RECT 42.445 4.115 42.695 5.125 ;
  LAYER M1 ;
        RECT 42.445 6.215 42.695 9.745 ;
  LAYER M1 ;
        RECT 42.445 9.995 42.695 11.005 ;
  LAYER M1 ;
        RECT 42.445 12.095 42.695 15.625 ;
  LAYER M1 ;
        RECT 42.445 15.875 42.695 16.885 ;
  LAYER M1 ;
        RECT 42.445 17.975 42.695 21.505 ;
  LAYER M1 ;
        RECT 42.445 21.755 42.695 22.765 ;
  LAYER M1 ;
        RECT 42.445 23.855 42.695 27.385 ;
  LAYER M1 ;
        RECT 42.445 27.635 42.695 28.645 ;
  LAYER M1 ;
        RECT 42.445 29.735 42.695 30.745 ;
  LAYER M1 ;
        RECT 42.875 0.335 43.125 3.865 ;
  LAYER M1 ;
        RECT 42.875 6.215 43.125 9.745 ;
  LAYER M1 ;
        RECT 42.875 12.095 43.125 15.625 ;
  LAYER M1 ;
        RECT 42.875 17.975 43.125 21.505 ;
  LAYER M1 ;
        RECT 42.875 23.855 43.125 27.385 ;
  LAYER M2 ;
        RECT 34.66 0.28 42.74 0.56 ;
  LAYER M2 ;
        RECT 34.66 4.48 42.74 4.76 ;
  LAYER M2 ;
        RECT 34.23 0.7 43.17 0.98 ;
  LAYER M2 ;
        RECT 34.66 6.16 42.74 6.44 ;
  LAYER M2 ;
        RECT 34.66 10.36 42.74 10.64 ;
  LAYER M2 ;
        RECT 34.23 6.58 43.17 6.86 ;
  LAYER M2 ;
        RECT 34.66 12.04 42.74 12.32 ;
  LAYER M2 ;
        RECT 34.66 16.24 42.74 16.52 ;
  LAYER M2 ;
        RECT 34.23 12.46 43.17 12.74 ;
  LAYER M2 ;
        RECT 34.66 17.92 42.74 18.2 ;
  LAYER M2 ;
        RECT 34.66 22.12 42.74 22.4 ;
  LAYER M2 ;
        RECT 34.23 18.34 43.17 18.62 ;
  LAYER M2 ;
        RECT 34.66 23.8 42.74 24.08 ;
  LAYER M2 ;
        RECT 34.66 28 42.74 28.28 ;
  LAYER M2 ;
        RECT 34.66 30.1 42.74 30.38 ;
  LAYER M2 ;
        RECT 34.23 24.22 43.17 24.5 ;
  LAYER M3 ;
        RECT 38.13 0.26 38.41 24.1 ;
  LAYER M3 ;
        RECT 38.56 4.46 38.84 28.3 ;
  LAYER M3 ;
        RECT 38.99 0.68 39.27 30.4 ;
  LAYER M1 ;
        RECT 21.805 27.215 22.055 30.745 ;
  LAYER M1 ;
        RECT 21.805 25.955 22.055 26.965 ;
  LAYER M1 ;
        RECT 21.805 21.335 22.055 24.865 ;
  LAYER M1 ;
        RECT 21.805 20.075 22.055 21.085 ;
  LAYER M1 ;
        RECT 21.805 17.975 22.055 18.985 ;
  LAYER M1 ;
        RECT 22.235 27.215 22.485 30.745 ;
  LAYER M1 ;
        RECT 22.235 21.335 22.485 24.865 ;
  LAYER M1 ;
        RECT 21.375 27.215 21.625 30.745 ;
  LAYER M1 ;
        RECT 21.375 21.335 21.625 24.865 ;
  LAYER M1 ;
        RECT 20.945 27.215 21.195 30.745 ;
  LAYER M1 ;
        RECT 20.945 25.955 21.195 26.965 ;
  LAYER M1 ;
        RECT 20.945 21.335 21.195 24.865 ;
  LAYER M1 ;
        RECT 20.945 20.075 21.195 21.085 ;
  LAYER M1 ;
        RECT 20.945 17.975 21.195 18.985 ;
  LAYER M1 ;
        RECT 20.515 27.215 20.765 30.745 ;
  LAYER M1 ;
        RECT 20.515 21.335 20.765 24.865 ;
  LAYER M1 ;
        RECT 20.085 27.215 20.335 30.745 ;
  LAYER M1 ;
        RECT 20.085 25.955 20.335 26.965 ;
  LAYER M1 ;
        RECT 20.085 21.335 20.335 24.865 ;
  LAYER M1 ;
        RECT 20.085 20.075 20.335 21.085 ;
  LAYER M1 ;
        RECT 20.085 17.975 20.335 18.985 ;
  LAYER M1 ;
        RECT 19.655 27.215 19.905 30.745 ;
  LAYER M1 ;
        RECT 19.655 21.335 19.905 24.865 ;
  LAYER M1 ;
        RECT 19.225 27.215 19.475 30.745 ;
  LAYER M1 ;
        RECT 19.225 25.955 19.475 26.965 ;
  LAYER M1 ;
        RECT 19.225 21.335 19.475 24.865 ;
  LAYER M1 ;
        RECT 19.225 20.075 19.475 21.085 ;
  LAYER M1 ;
        RECT 19.225 17.975 19.475 18.985 ;
  LAYER M1 ;
        RECT 18.795 27.215 19.045 30.745 ;
  LAYER M1 ;
        RECT 18.795 21.335 19.045 24.865 ;
  LAYER M1 ;
        RECT 18.365 27.215 18.615 30.745 ;
  LAYER M1 ;
        RECT 18.365 25.955 18.615 26.965 ;
  LAYER M1 ;
        RECT 18.365 21.335 18.615 24.865 ;
  LAYER M1 ;
        RECT 18.365 20.075 18.615 21.085 ;
  LAYER M1 ;
        RECT 18.365 17.975 18.615 18.985 ;
  LAYER M1 ;
        RECT 17.935 27.215 18.185 30.745 ;
  LAYER M1 ;
        RECT 17.935 21.335 18.185 24.865 ;
  LAYER M1 ;
        RECT 17.505 27.215 17.755 30.745 ;
  LAYER M1 ;
        RECT 17.505 25.955 17.755 26.965 ;
  LAYER M1 ;
        RECT 17.505 21.335 17.755 24.865 ;
  LAYER M1 ;
        RECT 17.505 20.075 17.755 21.085 ;
  LAYER M1 ;
        RECT 17.505 17.975 17.755 18.985 ;
  LAYER M1 ;
        RECT 17.075 27.215 17.325 30.745 ;
  LAYER M1 ;
        RECT 17.075 21.335 17.325 24.865 ;
  LAYER M1 ;
        RECT 16.645 27.215 16.895 30.745 ;
  LAYER M1 ;
        RECT 16.645 25.955 16.895 26.965 ;
  LAYER M1 ;
        RECT 16.645 21.335 16.895 24.865 ;
  LAYER M1 ;
        RECT 16.645 20.075 16.895 21.085 ;
  LAYER M1 ;
        RECT 16.645 17.975 16.895 18.985 ;
  LAYER M1 ;
        RECT 16.215 27.215 16.465 30.745 ;
  LAYER M1 ;
        RECT 16.215 21.335 16.465 24.865 ;
  LAYER M1 ;
        RECT 15.785 27.215 16.035 30.745 ;
  LAYER M1 ;
        RECT 15.785 25.955 16.035 26.965 ;
  LAYER M1 ;
        RECT 15.785 21.335 16.035 24.865 ;
  LAYER M1 ;
        RECT 15.785 20.075 16.035 21.085 ;
  LAYER M1 ;
        RECT 15.785 17.975 16.035 18.985 ;
  LAYER M1 ;
        RECT 15.355 27.215 15.605 30.745 ;
  LAYER M1 ;
        RECT 15.355 21.335 15.605 24.865 ;
  LAYER M1 ;
        RECT 14.925 27.215 15.175 30.745 ;
  LAYER M1 ;
        RECT 14.925 25.955 15.175 26.965 ;
  LAYER M1 ;
        RECT 14.925 21.335 15.175 24.865 ;
  LAYER M1 ;
        RECT 14.925 20.075 15.175 21.085 ;
  LAYER M1 ;
        RECT 14.925 17.975 15.175 18.985 ;
  LAYER M1 ;
        RECT 14.495 27.215 14.745 30.745 ;
  LAYER M1 ;
        RECT 14.495 21.335 14.745 24.865 ;
  LAYER M1 ;
        RECT 14.065 27.215 14.315 30.745 ;
  LAYER M1 ;
        RECT 14.065 25.955 14.315 26.965 ;
  LAYER M1 ;
        RECT 14.065 21.335 14.315 24.865 ;
  LAYER M1 ;
        RECT 14.065 20.075 14.315 21.085 ;
  LAYER M1 ;
        RECT 14.065 17.975 14.315 18.985 ;
  LAYER M1 ;
        RECT 13.635 27.215 13.885 30.745 ;
  LAYER M1 ;
        RECT 13.635 21.335 13.885 24.865 ;
  LAYER M1 ;
        RECT 13.205 27.215 13.455 30.745 ;
  LAYER M1 ;
        RECT 13.205 25.955 13.455 26.965 ;
  LAYER M1 ;
        RECT 13.205 21.335 13.455 24.865 ;
  LAYER M1 ;
        RECT 13.205 20.075 13.455 21.085 ;
  LAYER M1 ;
        RECT 13.205 17.975 13.455 18.985 ;
  LAYER M1 ;
        RECT 12.775 27.215 13.025 30.745 ;
  LAYER M1 ;
        RECT 12.775 21.335 13.025 24.865 ;
  LAYER M1 ;
        RECT 12.345 27.215 12.595 30.745 ;
  LAYER M1 ;
        RECT 12.345 25.955 12.595 26.965 ;
  LAYER M1 ;
        RECT 12.345 21.335 12.595 24.865 ;
  LAYER M1 ;
        RECT 12.345 20.075 12.595 21.085 ;
  LAYER M1 ;
        RECT 12.345 17.975 12.595 18.985 ;
  LAYER M1 ;
        RECT 11.915 27.215 12.165 30.745 ;
  LAYER M1 ;
        RECT 11.915 21.335 12.165 24.865 ;
  LAYER M1 ;
        RECT 11.485 27.215 11.735 30.745 ;
  LAYER M1 ;
        RECT 11.485 25.955 11.735 26.965 ;
  LAYER M1 ;
        RECT 11.485 21.335 11.735 24.865 ;
  LAYER M1 ;
        RECT 11.485 20.075 11.735 21.085 ;
  LAYER M1 ;
        RECT 11.485 17.975 11.735 18.985 ;
  LAYER M1 ;
        RECT 11.055 27.215 11.305 30.745 ;
  LAYER M1 ;
        RECT 11.055 21.335 11.305 24.865 ;
  LAYER M1 ;
        RECT 10.625 27.215 10.875 30.745 ;
  LAYER M1 ;
        RECT 10.625 25.955 10.875 26.965 ;
  LAYER M1 ;
        RECT 10.625 21.335 10.875 24.865 ;
  LAYER M1 ;
        RECT 10.625 20.075 10.875 21.085 ;
  LAYER M1 ;
        RECT 10.625 17.975 10.875 18.985 ;
  LAYER M1 ;
        RECT 10.195 27.215 10.445 30.745 ;
  LAYER M1 ;
        RECT 10.195 21.335 10.445 24.865 ;
  LAYER M1 ;
        RECT 9.765 27.215 10.015 30.745 ;
  LAYER M1 ;
        RECT 9.765 25.955 10.015 26.965 ;
  LAYER M1 ;
        RECT 9.765 21.335 10.015 24.865 ;
  LAYER M1 ;
        RECT 9.765 20.075 10.015 21.085 ;
  LAYER M1 ;
        RECT 9.765 17.975 10.015 18.985 ;
  LAYER M1 ;
        RECT 9.335 27.215 9.585 30.745 ;
  LAYER M1 ;
        RECT 9.335 21.335 9.585 24.865 ;
  LAYER M1 ;
        RECT 8.905 27.215 9.155 30.745 ;
  LAYER M1 ;
        RECT 8.905 25.955 9.155 26.965 ;
  LAYER M1 ;
        RECT 8.905 21.335 9.155 24.865 ;
  LAYER M1 ;
        RECT 8.905 20.075 9.155 21.085 ;
  LAYER M1 ;
        RECT 8.905 17.975 9.155 18.985 ;
  LAYER M1 ;
        RECT 8.475 27.215 8.725 30.745 ;
  LAYER M1 ;
        RECT 8.475 21.335 8.725 24.865 ;
  LAYER M1 ;
        RECT 8.045 27.215 8.295 30.745 ;
  LAYER M1 ;
        RECT 8.045 25.955 8.295 26.965 ;
  LAYER M1 ;
        RECT 8.045 21.335 8.295 24.865 ;
  LAYER M1 ;
        RECT 8.045 20.075 8.295 21.085 ;
  LAYER M1 ;
        RECT 8.045 17.975 8.295 18.985 ;
  LAYER M1 ;
        RECT 7.615 27.215 7.865 30.745 ;
  LAYER M1 ;
        RECT 7.615 21.335 7.865 24.865 ;
  LAYER M1 ;
        RECT 7.185 27.215 7.435 30.745 ;
  LAYER M1 ;
        RECT 7.185 25.955 7.435 26.965 ;
  LAYER M1 ;
        RECT 7.185 21.335 7.435 24.865 ;
  LAYER M1 ;
        RECT 7.185 20.075 7.435 21.085 ;
  LAYER M1 ;
        RECT 7.185 17.975 7.435 18.985 ;
  LAYER M1 ;
        RECT 6.755 27.215 7.005 30.745 ;
  LAYER M1 ;
        RECT 6.755 21.335 7.005 24.865 ;
  LAYER M2 ;
        RECT 7.14 30.52 22.1 30.8 ;
  LAYER M2 ;
        RECT 7.14 26.32 22.1 26.6 ;
  LAYER M2 ;
        RECT 6.71 30.1 22.53 30.38 ;
  LAYER M2 ;
        RECT 7.14 24.64 22.1 24.92 ;
  LAYER M2 ;
        RECT 7.14 20.44 22.1 20.72 ;
  LAYER M2 ;
        RECT 7.14 18.34 22.1 18.62 ;
  LAYER M2 ;
        RECT 6.71 24.22 22.53 24.5 ;
  LAYER M3 ;
        RECT 14.91 24.62 15.19 30.82 ;
  LAYER M3 ;
        RECT 14.48 20.42 14.76 26.62 ;
  LAYER M3 ;
        RECT 14.05 18.32 14.33 30.4 ;
  LAYER M1 ;
        RECT 45.025 27.215 45.275 30.745 ;
  LAYER M1 ;
        RECT 45.025 25.955 45.275 26.965 ;
  LAYER M1 ;
        RECT 45.025 21.335 45.275 24.865 ;
  LAYER M1 ;
        RECT 45.025 20.075 45.275 21.085 ;
  LAYER M1 ;
        RECT 45.025 17.975 45.275 18.985 ;
  LAYER M1 ;
        RECT 44.595 27.215 44.845 30.745 ;
  LAYER M1 ;
        RECT 44.595 21.335 44.845 24.865 ;
  LAYER M1 ;
        RECT 45.455 27.215 45.705 30.745 ;
  LAYER M1 ;
        RECT 45.455 21.335 45.705 24.865 ;
  LAYER M1 ;
        RECT 45.885 27.215 46.135 30.745 ;
  LAYER M1 ;
        RECT 45.885 25.955 46.135 26.965 ;
  LAYER M1 ;
        RECT 45.885 21.335 46.135 24.865 ;
  LAYER M1 ;
        RECT 45.885 20.075 46.135 21.085 ;
  LAYER M1 ;
        RECT 45.885 17.975 46.135 18.985 ;
  LAYER M1 ;
        RECT 46.315 27.215 46.565 30.745 ;
  LAYER M1 ;
        RECT 46.315 21.335 46.565 24.865 ;
  LAYER M1 ;
        RECT 46.745 27.215 46.995 30.745 ;
  LAYER M1 ;
        RECT 46.745 25.955 46.995 26.965 ;
  LAYER M1 ;
        RECT 46.745 21.335 46.995 24.865 ;
  LAYER M1 ;
        RECT 46.745 20.075 46.995 21.085 ;
  LAYER M1 ;
        RECT 46.745 17.975 46.995 18.985 ;
  LAYER M1 ;
        RECT 47.175 27.215 47.425 30.745 ;
  LAYER M1 ;
        RECT 47.175 21.335 47.425 24.865 ;
  LAYER M1 ;
        RECT 47.605 27.215 47.855 30.745 ;
  LAYER M1 ;
        RECT 47.605 25.955 47.855 26.965 ;
  LAYER M1 ;
        RECT 47.605 21.335 47.855 24.865 ;
  LAYER M1 ;
        RECT 47.605 20.075 47.855 21.085 ;
  LAYER M1 ;
        RECT 47.605 17.975 47.855 18.985 ;
  LAYER M1 ;
        RECT 48.035 27.215 48.285 30.745 ;
  LAYER M1 ;
        RECT 48.035 21.335 48.285 24.865 ;
  LAYER M1 ;
        RECT 48.465 27.215 48.715 30.745 ;
  LAYER M1 ;
        RECT 48.465 25.955 48.715 26.965 ;
  LAYER M1 ;
        RECT 48.465 21.335 48.715 24.865 ;
  LAYER M1 ;
        RECT 48.465 20.075 48.715 21.085 ;
  LAYER M1 ;
        RECT 48.465 17.975 48.715 18.985 ;
  LAYER M1 ;
        RECT 48.895 27.215 49.145 30.745 ;
  LAYER M1 ;
        RECT 48.895 21.335 49.145 24.865 ;
  LAYER M1 ;
        RECT 49.325 27.215 49.575 30.745 ;
  LAYER M1 ;
        RECT 49.325 25.955 49.575 26.965 ;
  LAYER M1 ;
        RECT 49.325 21.335 49.575 24.865 ;
  LAYER M1 ;
        RECT 49.325 20.075 49.575 21.085 ;
  LAYER M1 ;
        RECT 49.325 17.975 49.575 18.985 ;
  LAYER M1 ;
        RECT 49.755 27.215 50.005 30.745 ;
  LAYER M1 ;
        RECT 49.755 21.335 50.005 24.865 ;
  LAYER M1 ;
        RECT 50.185 27.215 50.435 30.745 ;
  LAYER M1 ;
        RECT 50.185 25.955 50.435 26.965 ;
  LAYER M1 ;
        RECT 50.185 21.335 50.435 24.865 ;
  LAYER M1 ;
        RECT 50.185 20.075 50.435 21.085 ;
  LAYER M1 ;
        RECT 50.185 17.975 50.435 18.985 ;
  LAYER M1 ;
        RECT 50.615 27.215 50.865 30.745 ;
  LAYER M1 ;
        RECT 50.615 21.335 50.865 24.865 ;
  LAYER M1 ;
        RECT 51.045 27.215 51.295 30.745 ;
  LAYER M1 ;
        RECT 51.045 25.955 51.295 26.965 ;
  LAYER M1 ;
        RECT 51.045 21.335 51.295 24.865 ;
  LAYER M1 ;
        RECT 51.045 20.075 51.295 21.085 ;
  LAYER M1 ;
        RECT 51.045 17.975 51.295 18.985 ;
  LAYER M1 ;
        RECT 51.475 27.215 51.725 30.745 ;
  LAYER M1 ;
        RECT 51.475 21.335 51.725 24.865 ;
  LAYER M1 ;
        RECT 51.905 27.215 52.155 30.745 ;
  LAYER M1 ;
        RECT 51.905 25.955 52.155 26.965 ;
  LAYER M1 ;
        RECT 51.905 21.335 52.155 24.865 ;
  LAYER M1 ;
        RECT 51.905 20.075 52.155 21.085 ;
  LAYER M1 ;
        RECT 51.905 17.975 52.155 18.985 ;
  LAYER M1 ;
        RECT 52.335 27.215 52.585 30.745 ;
  LAYER M1 ;
        RECT 52.335 21.335 52.585 24.865 ;
  LAYER M1 ;
        RECT 52.765 27.215 53.015 30.745 ;
  LAYER M1 ;
        RECT 52.765 25.955 53.015 26.965 ;
  LAYER M1 ;
        RECT 52.765 21.335 53.015 24.865 ;
  LAYER M1 ;
        RECT 52.765 20.075 53.015 21.085 ;
  LAYER M1 ;
        RECT 52.765 17.975 53.015 18.985 ;
  LAYER M1 ;
        RECT 53.195 27.215 53.445 30.745 ;
  LAYER M1 ;
        RECT 53.195 21.335 53.445 24.865 ;
  LAYER M1 ;
        RECT 53.625 27.215 53.875 30.745 ;
  LAYER M1 ;
        RECT 53.625 25.955 53.875 26.965 ;
  LAYER M1 ;
        RECT 53.625 21.335 53.875 24.865 ;
  LAYER M1 ;
        RECT 53.625 20.075 53.875 21.085 ;
  LAYER M1 ;
        RECT 53.625 17.975 53.875 18.985 ;
  LAYER M1 ;
        RECT 54.055 27.215 54.305 30.745 ;
  LAYER M1 ;
        RECT 54.055 21.335 54.305 24.865 ;
  LAYER M1 ;
        RECT 54.485 27.215 54.735 30.745 ;
  LAYER M1 ;
        RECT 54.485 25.955 54.735 26.965 ;
  LAYER M1 ;
        RECT 54.485 21.335 54.735 24.865 ;
  LAYER M1 ;
        RECT 54.485 20.075 54.735 21.085 ;
  LAYER M1 ;
        RECT 54.485 17.975 54.735 18.985 ;
  LAYER M1 ;
        RECT 54.915 27.215 55.165 30.745 ;
  LAYER M1 ;
        RECT 54.915 21.335 55.165 24.865 ;
  LAYER M1 ;
        RECT 55.345 27.215 55.595 30.745 ;
  LAYER M1 ;
        RECT 55.345 25.955 55.595 26.965 ;
  LAYER M1 ;
        RECT 55.345 21.335 55.595 24.865 ;
  LAYER M1 ;
        RECT 55.345 20.075 55.595 21.085 ;
  LAYER M1 ;
        RECT 55.345 17.975 55.595 18.985 ;
  LAYER M1 ;
        RECT 55.775 27.215 56.025 30.745 ;
  LAYER M1 ;
        RECT 55.775 21.335 56.025 24.865 ;
  LAYER M1 ;
        RECT 56.205 27.215 56.455 30.745 ;
  LAYER M1 ;
        RECT 56.205 25.955 56.455 26.965 ;
  LAYER M1 ;
        RECT 56.205 21.335 56.455 24.865 ;
  LAYER M1 ;
        RECT 56.205 20.075 56.455 21.085 ;
  LAYER M1 ;
        RECT 56.205 17.975 56.455 18.985 ;
  LAYER M1 ;
        RECT 56.635 27.215 56.885 30.745 ;
  LAYER M1 ;
        RECT 56.635 21.335 56.885 24.865 ;
  LAYER M1 ;
        RECT 57.065 27.215 57.315 30.745 ;
  LAYER M1 ;
        RECT 57.065 25.955 57.315 26.965 ;
  LAYER M1 ;
        RECT 57.065 21.335 57.315 24.865 ;
  LAYER M1 ;
        RECT 57.065 20.075 57.315 21.085 ;
  LAYER M1 ;
        RECT 57.065 17.975 57.315 18.985 ;
  LAYER M1 ;
        RECT 57.495 27.215 57.745 30.745 ;
  LAYER M1 ;
        RECT 57.495 21.335 57.745 24.865 ;
  LAYER M1 ;
        RECT 57.925 27.215 58.175 30.745 ;
  LAYER M1 ;
        RECT 57.925 25.955 58.175 26.965 ;
  LAYER M1 ;
        RECT 57.925 21.335 58.175 24.865 ;
  LAYER M1 ;
        RECT 57.925 20.075 58.175 21.085 ;
  LAYER M1 ;
        RECT 57.925 17.975 58.175 18.985 ;
  LAYER M1 ;
        RECT 58.355 27.215 58.605 30.745 ;
  LAYER M1 ;
        RECT 58.355 21.335 58.605 24.865 ;
  LAYER M1 ;
        RECT 58.785 27.215 59.035 30.745 ;
  LAYER M1 ;
        RECT 58.785 25.955 59.035 26.965 ;
  LAYER M1 ;
        RECT 58.785 21.335 59.035 24.865 ;
  LAYER M1 ;
        RECT 58.785 20.075 59.035 21.085 ;
  LAYER M1 ;
        RECT 58.785 17.975 59.035 18.985 ;
  LAYER M1 ;
        RECT 59.215 27.215 59.465 30.745 ;
  LAYER M1 ;
        RECT 59.215 21.335 59.465 24.865 ;
  LAYER M1 ;
        RECT 59.645 27.215 59.895 30.745 ;
  LAYER M1 ;
        RECT 59.645 25.955 59.895 26.965 ;
  LAYER M1 ;
        RECT 59.645 21.335 59.895 24.865 ;
  LAYER M1 ;
        RECT 59.645 20.075 59.895 21.085 ;
  LAYER M1 ;
        RECT 59.645 17.975 59.895 18.985 ;
  LAYER M1 ;
        RECT 60.075 27.215 60.325 30.745 ;
  LAYER M1 ;
        RECT 60.075 21.335 60.325 24.865 ;
  LAYER M2 ;
        RECT 44.98 30.52 59.94 30.8 ;
  LAYER M2 ;
        RECT 44.98 26.32 59.94 26.6 ;
  LAYER M2 ;
        RECT 44.55 30.1 60.37 30.38 ;
  LAYER M2 ;
        RECT 44.98 24.64 59.94 24.92 ;
  LAYER M2 ;
        RECT 44.98 20.44 59.94 20.72 ;
  LAYER M2 ;
        RECT 44.98 18.34 59.94 18.62 ;
  LAYER M2 ;
        RECT 44.55 24.22 60.37 24.5 ;
  LAYER M3 ;
        RECT 51.89 24.62 52.17 30.82 ;
  LAYER M3 ;
        RECT 52.32 20.42 52.6 26.62 ;
  LAYER M3 ;
        RECT 52.75 18.32 53.03 30.4 ;
  LAYER M1 ;
        RECT 21.805 12.095 22.055 15.625 ;
  LAYER M1 ;
        RECT 21.805 10.835 22.055 11.845 ;
  LAYER M1 ;
        RECT 21.805 8.735 22.055 9.745 ;
  LAYER M1 ;
        RECT 22.235 12.095 22.485 15.625 ;
  LAYER M1 ;
        RECT 21.375 12.095 21.625 15.625 ;
  LAYER M1 ;
        RECT 20.945 12.095 21.195 15.625 ;
  LAYER M1 ;
        RECT 20.945 10.835 21.195 11.845 ;
  LAYER M1 ;
        RECT 20.945 8.735 21.195 9.745 ;
  LAYER M1 ;
        RECT 20.515 12.095 20.765 15.625 ;
  LAYER M1 ;
        RECT 20.085 12.095 20.335 15.625 ;
  LAYER M1 ;
        RECT 20.085 10.835 20.335 11.845 ;
  LAYER M1 ;
        RECT 20.085 8.735 20.335 9.745 ;
  LAYER M1 ;
        RECT 19.655 12.095 19.905 15.625 ;
  LAYER M1 ;
        RECT 19.225 12.095 19.475 15.625 ;
  LAYER M1 ;
        RECT 19.225 10.835 19.475 11.845 ;
  LAYER M1 ;
        RECT 19.225 8.735 19.475 9.745 ;
  LAYER M1 ;
        RECT 18.795 12.095 19.045 15.625 ;
  LAYER M1 ;
        RECT 18.365 12.095 18.615 15.625 ;
  LAYER M1 ;
        RECT 18.365 10.835 18.615 11.845 ;
  LAYER M1 ;
        RECT 18.365 8.735 18.615 9.745 ;
  LAYER M1 ;
        RECT 17.935 12.095 18.185 15.625 ;
  LAYER M1 ;
        RECT 17.505 12.095 17.755 15.625 ;
  LAYER M1 ;
        RECT 17.505 10.835 17.755 11.845 ;
  LAYER M1 ;
        RECT 17.505 8.735 17.755 9.745 ;
  LAYER M1 ;
        RECT 17.075 12.095 17.325 15.625 ;
  LAYER M1 ;
        RECT 16.645 12.095 16.895 15.625 ;
  LAYER M1 ;
        RECT 16.645 10.835 16.895 11.845 ;
  LAYER M1 ;
        RECT 16.645 8.735 16.895 9.745 ;
  LAYER M1 ;
        RECT 16.215 12.095 16.465 15.625 ;
  LAYER M1 ;
        RECT 15.785 12.095 16.035 15.625 ;
  LAYER M1 ;
        RECT 15.785 10.835 16.035 11.845 ;
  LAYER M1 ;
        RECT 15.785 8.735 16.035 9.745 ;
  LAYER M1 ;
        RECT 15.355 12.095 15.605 15.625 ;
  LAYER M1 ;
        RECT 14.925 12.095 15.175 15.625 ;
  LAYER M1 ;
        RECT 14.925 10.835 15.175 11.845 ;
  LAYER M1 ;
        RECT 14.925 8.735 15.175 9.745 ;
  LAYER M1 ;
        RECT 14.495 12.095 14.745 15.625 ;
  LAYER M1 ;
        RECT 14.065 12.095 14.315 15.625 ;
  LAYER M1 ;
        RECT 14.065 10.835 14.315 11.845 ;
  LAYER M1 ;
        RECT 14.065 8.735 14.315 9.745 ;
  LAYER M1 ;
        RECT 13.635 12.095 13.885 15.625 ;
  LAYER M1 ;
        RECT 13.205 12.095 13.455 15.625 ;
  LAYER M1 ;
        RECT 13.205 10.835 13.455 11.845 ;
  LAYER M1 ;
        RECT 13.205 8.735 13.455 9.745 ;
  LAYER M1 ;
        RECT 12.775 12.095 13.025 15.625 ;
  LAYER M1 ;
        RECT 12.345 12.095 12.595 15.625 ;
  LAYER M1 ;
        RECT 12.345 10.835 12.595 11.845 ;
  LAYER M1 ;
        RECT 12.345 8.735 12.595 9.745 ;
  LAYER M1 ;
        RECT 11.915 12.095 12.165 15.625 ;
  LAYER M1 ;
        RECT 11.485 12.095 11.735 15.625 ;
  LAYER M1 ;
        RECT 11.485 10.835 11.735 11.845 ;
  LAYER M1 ;
        RECT 11.485 8.735 11.735 9.745 ;
  LAYER M1 ;
        RECT 11.055 12.095 11.305 15.625 ;
  LAYER M1 ;
        RECT 10.625 12.095 10.875 15.625 ;
  LAYER M1 ;
        RECT 10.625 10.835 10.875 11.845 ;
  LAYER M1 ;
        RECT 10.625 8.735 10.875 9.745 ;
  LAYER M1 ;
        RECT 10.195 12.095 10.445 15.625 ;
  LAYER M1 ;
        RECT 9.765 12.095 10.015 15.625 ;
  LAYER M1 ;
        RECT 9.765 10.835 10.015 11.845 ;
  LAYER M1 ;
        RECT 9.765 8.735 10.015 9.745 ;
  LAYER M1 ;
        RECT 9.335 12.095 9.585 15.625 ;
  LAYER M1 ;
        RECT 8.905 12.095 9.155 15.625 ;
  LAYER M1 ;
        RECT 8.905 10.835 9.155 11.845 ;
  LAYER M1 ;
        RECT 8.905 8.735 9.155 9.745 ;
  LAYER M1 ;
        RECT 8.475 12.095 8.725 15.625 ;
  LAYER M1 ;
        RECT 8.045 12.095 8.295 15.625 ;
  LAYER M1 ;
        RECT 8.045 10.835 8.295 11.845 ;
  LAYER M1 ;
        RECT 8.045 8.735 8.295 9.745 ;
  LAYER M1 ;
        RECT 7.615 12.095 7.865 15.625 ;
  LAYER M1 ;
        RECT 7.185 12.095 7.435 15.625 ;
  LAYER M1 ;
        RECT 7.185 10.835 7.435 11.845 ;
  LAYER M1 ;
        RECT 7.185 8.735 7.435 9.745 ;
  LAYER M1 ;
        RECT 6.755 12.095 7.005 15.625 ;
  LAYER M1 ;
        RECT 6.325 12.095 6.575 15.625 ;
  LAYER M1 ;
        RECT 6.325 10.835 6.575 11.845 ;
  LAYER M1 ;
        RECT 6.325 8.735 6.575 9.745 ;
  LAYER M1 ;
        RECT 5.895 12.095 6.145 15.625 ;
  LAYER M1 ;
        RECT 5.465 12.095 5.715 15.625 ;
  LAYER M1 ;
        RECT 5.465 10.835 5.715 11.845 ;
  LAYER M1 ;
        RECT 5.465 8.735 5.715 9.745 ;
  LAYER M1 ;
        RECT 5.035 12.095 5.285 15.625 ;
  LAYER M1 ;
        RECT 4.605 12.095 4.855 15.625 ;
  LAYER M1 ;
        RECT 4.605 10.835 4.855 11.845 ;
  LAYER M1 ;
        RECT 4.605 8.735 4.855 9.745 ;
  LAYER M1 ;
        RECT 4.175 12.095 4.425 15.625 ;
  LAYER M1 ;
        RECT 3.745 12.095 3.995 15.625 ;
  LAYER M1 ;
        RECT 3.745 10.835 3.995 11.845 ;
  LAYER M1 ;
        RECT 3.745 8.735 3.995 9.745 ;
  LAYER M1 ;
        RECT 3.315 12.095 3.565 15.625 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 15.625 ;
  LAYER M1 ;
        RECT 2.885 10.835 3.135 11.845 ;
  LAYER M1 ;
        RECT 2.885 8.735 3.135 9.745 ;
  LAYER M1 ;
        RECT 2.455 12.095 2.705 15.625 ;
  LAYER M1 ;
        RECT 2.025 12.095 2.275 15.625 ;
  LAYER M1 ;
        RECT 2.025 10.835 2.275 11.845 ;
  LAYER M1 ;
        RECT 2.025 8.735 2.275 9.745 ;
  LAYER M1 ;
        RECT 1.595 12.095 1.845 15.625 ;
  LAYER M1 ;
        RECT 1.165 12.095 1.415 15.625 ;
  LAYER M1 ;
        RECT 1.165 10.835 1.415 11.845 ;
  LAYER M1 ;
        RECT 1.165 8.735 1.415 9.745 ;
  LAYER M1 ;
        RECT 0.735 12.095 0.985 15.625 ;
  LAYER M2 ;
        RECT 1.12 9.1 22.1 9.38 ;
  LAYER M2 ;
        RECT 1.12 15.4 22.1 15.68 ;
  LAYER M2 ;
        RECT 1.12 11.2 22.1 11.48 ;
  LAYER M2 ;
        RECT 0.69 14.98 22.53 15.26 ;
  LAYER M1 ;
        RECT 45.025 12.095 45.275 15.625 ;
  LAYER M1 ;
        RECT 45.025 10.835 45.275 11.845 ;
  LAYER M1 ;
        RECT 45.025 8.735 45.275 9.745 ;
  LAYER M1 ;
        RECT 44.595 12.095 44.845 15.625 ;
  LAYER M1 ;
        RECT 45.455 12.095 45.705 15.625 ;
  LAYER M1 ;
        RECT 45.885 12.095 46.135 15.625 ;
  LAYER M1 ;
        RECT 45.885 10.835 46.135 11.845 ;
  LAYER M1 ;
        RECT 45.885 8.735 46.135 9.745 ;
  LAYER M1 ;
        RECT 46.315 12.095 46.565 15.625 ;
  LAYER M1 ;
        RECT 46.745 12.095 46.995 15.625 ;
  LAYER M1 ;
        RECT 46.745 10.835 46.995 11.845 ;
  LAYER M1 ;
        RECT 46.745 8.735 46.995 9.745 ;
  LAYER M1 ;
        RECT 47.175 12.095 47.425 15.625 ;
  LAYER M1 ;
        RECT 47.605 12.095 47.855 15.625 ;
  LAYER M1 ;
        RECT 47.605 10.835 47.855 11.845 ;
  LAYER M1 ;
        RECT 47.605 8.735 47.855 9.745 ;
  LAYER M1 ;
        RECT 48.035 12.095 48.285 15.625 ;
  LAYER M1 ;
        RECT 48.465 12.095 48.715 15.625 ;
  LAYER M1 ;
        RECT 48.465 10.835 48.715 11.845 ;
  LAYER M1 ;
        RECT 48.465 8.735 48.715 9.745 ;
  LAYER M1 ;
        RECT 48.895 12.095 49.145 15.625 ;
  LAYER M1 ;
        RECT 49.325 12.095 49.575 15.625 ;
  LAYER M1 ;
        RECT 49.325 10.835 49.575 11.845 ;
  LAYER M1 ;
        RECT 49.325 8.735 49.575 9.745 ;
  LAYER M1 ;
        RECT 49.755 12.095 50.005 15.625 ;
  LAYER M1 ;
        RECT 50.185 12.095 50.435 15.625 ;
  LAYER M1 ;
        RECT 50.185 10.835 50.435 11.845 ;
  LAYER M1 ;
        RECT 50.185 8.735 50.435 9.745 ;
  LAYER M1 ;
        RECT 50.615 12.095 50.865 15.625 ;
  LAYER M1 ;
        RECT 51.045 12.095 51.295 15.625 ;
  LAYER M1 ;
        RECT 51.045 10.835 51.295 11.845 ;
  LAYER M1 ;
        RECT 51.045 8.735 51.295 9.745 ;
  LAYER M1 ;
        RECT 51.475 12.095 51.725 15.625 ;
  LAYER M1 ;
        RECT 51.905 12.095 52.155 15.625 ;
  LAYER M1 ;
        RECT 51.905 10.835 52.155 11.845 ;
  LAYER M1 ;
        RECT 51.905 8.735 52.155 9.745 ;
  LAYER M1 ;
        RECT 52.335 12.095 52.585 15.625 ;
  LAYER M1 ;
        RECT 52.765 12.095 53.015 15.625 ;
  LAYER M1 ;
        RECT 52.765 10.835 53.015 11.845 ;
  LAYER M1 ;
        RECT 52.765 8.735 53.015 9.745 ;
  LAYER M1 ;
        RECT 53.195 12.095 53.445 15.625 ;
  LAYER M1 ;
        RECT 53.625 12.095 53.875 15.625 ;
  LAYER M1 ;
        RECT 53.625 10.835 53.875 11.845 ;
  LAYER M1 ;
        RECT 53.625 8.735 53.875 9.745 ;
  LAYER M1 ;
        RECT 54.055 12.095 54.305 15.625 ;
  LAYER M1 ;
        RECT 54.485 12.095 54.735 15.625 ;
  LAYER M1 ;
        RECT 54.485 10.835 54.735 11.845 ;
  LAYER M1 ;
        RECT 54.485 8.735 54.735 9.745 ;
  LAYER M1 ;
        RECT 54.915 12.095 55.165 15.625 ;
  LAYER M1 ;
        RECT 55.345 12.095 55.595 15.625 ;
  LAYER M1 ;
        RECT 55.345 10.835 55.595 11.845 ;
  LAYER M1 ;
        RECT 55.345 8.735 55.595 9.745 ;
  LAYER M1 ;
        RECT 55.775 12.095 56.025 15.625 ;
  LAYER M1 ;
        RECT 56.205 12.095 56.455 15.625 ;
  LAYER M1 ;
        RECT 56.205 10.835 56.455 11.845 ;
  LAYER M1 ;
        RECT 56.205 8.735 56.455 9.745 ;
  LAYER M1 ;
        RECT 56.635 12.095 56.885 15.625 ;
  LAYER M1 ;
        RECT 57.065 12.095 57.315 15.625 ;
  LAYER M1 ;
        RECT 57.065 10.835 57.315 11.845 ;
  LAYER M1 ;
        RECT 57.065 8.735 57.315 9.745 ;
  LAYER M1 ;
        RECT 57.495 12.095 57.745 15.625 ;
  LAYER M1 ;
        RECT 57.925 12.095 58.175 15.625 ;
  LAYER M1 ;
        RECT 57.925 10.835 58.175 11.845 ;
  LAYER M1 ;
        RECT 57.925 8.735 58.175 9.745 ;
  LAYER M1 ;
        RECT 58.355 12.095 58.605 15.625 ;
  LAYER M1 ;
        RECT 58.785 12.095 59.035 15.625 ;
  LAYER M1 ;
        RECT 58.785 10.835 59.035 11.845 ;
  LAYER M1 ;
        RECT 58.785 8.735 59.035 9.745 ;
  LAYER M1 ;
        RECT 59.215 12.095 59.465 15.625 ;
  LAYER M1 ;
        RECT 59.645 12.095 59.895 15.625 ;
  LAYER M1 ;
        RECT 59.645 10.835 59.895 11.845 ;
  LAYER M1 ;
        RECT 59.645 8.735 59.895 9.745 ;
  LAYER M1 ;
        RECT 60.075 12.095 60.325 15.625 ;
  LAYER M1 ;
        RECT 60.505 12.095 60.755 15.625 ;
  LAYER M1 ;
        RECT 60.505 10.835 60.755 11.845 ;
  LAYER M1 ;
        RECT 60.505 8.735 60.755 9.745 ;
  LAYER M1 ;
        RECT 60.935 12.095 61.185 15.625 ;
  LAYER M1 ;
        RECT 61.365 12.095 61.615 15.625 ;
  LAYER M1 ;
        RECT 61.365 10.835 61.615 11.845 ;
  LAYER M1 ;
        RECT 61.365 8.735 61.615 9.745 ;
  LAYER M1 ;
        RECT 61.795 12.095 62.045 15.625 ;
  LAYER M1 ;
        RECT 62.225 12.095 62.475 15.625 ;
  LAYER M1 ;
        RECT 62.225 10.835 62.475 11.845 ;
  LAYER M1 ;
        RECT 62.225 8.735 62.475 9.745 ;
  LAYER M1 ;
        RECT 62.655 12.095 62.905 15.625 ;
  LAYER M1 ;
        RECT 63.085 12.095 63.335 15.625 ;
  LAYER M1 ;
        RECT 63.085 10.835 63.335 11.845 ;
  LAYER M1 ;
        RECT 63.085 8.735 63.335 9.745 ;
  LAYER M1 ;
        RECT 63.515 12.095 63.765 15.625 ;
  LAYER M1 ;
        RECT 63.945 12.095 64.195 15.625 ;
  LAYER M1 ;
        RECT 63.945 10.835 64.195 11.845 ;
  LAYER M1 ;
        RECT 63.945 8.735 64.195 9.745 ;
  LAYER M1 ;
        RECT 64.375 12.095 64.625 15.625 ;
  LAYER M1 ;
        RECT 64.805 12.095 65.055 15.625 ;
  LAYER M1 ;
        RECT 64.805 10.835 65.055 11.845 ;
  LAYER M1 ;
        RECT 64.805 8.735 65.055 9.745 ;
  LAYER M1 ;
        RECT 65.235 12.095 65.485 15.625 ;
  LAYER M1 ;
        RECT 65.665 12.095 65.915 15.625 ;
  LAYER M1 ;
        RECT 65.665 10.835 65.915 11.845 ;
  LAYER M1 ;
        RECT 65.665 8.735 65.915 9.745 ;
  LAYER M1 ;
        RECT 66.095 12.095 66.345 15.625 ;
  LAYER M2 ;
        RECT 44.98 9.1 65.96 9.38 ;
  LAYER M2 ;
        RECT 44.98 15.4 65.96 15.68 ;
  LAYER M2 ;
        RECT 44.98 11.2 65.96 11.48 ;
  LAYER M2 ;
        RECT 44.55 14.98 66.39 15.26 ;
  END 
END CURRENT_MIRROR_OTA
