MACRO DCL_NMOS_S_38019457_X1_Y50
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_S_38019457_X1_Y50 0 0 ;
  SIZE 2580 BY 295680 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 260 1430 292900 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 295000 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 62665 ;
    LAYER M1 ;
      RECT 1165 62915 1415 63925 ;
    LAYER M1 ;
      RECT 1165 65015 1415 68545 ;
    LAYER M1 ;
      RECT 1165 68795 1415 69805 ;
    LAYER M1 ;
      RECT 1165 70895 1415 74425 ;
    LAYER M1 ;
      RECT 1165 74675 1415 75685 ;
    LAYER M1 ;
      RECT 1165 76775 1415 80305 ;
    LAYER M1 ;
      RECT 1165 80555 1415 81565 ;
    LAYER M1 ;
      RECT 1165 82655 1415 86185 ;
    LAYER M1 ;
      RECT 1165 86435 1415 87445 ;
    LAYER M1 ;
      RECT 1165 88535 1415 92065 ;
    LAYER M1 ;
      RECT 1165 92315 1415 93325 ;
    LAYER M1 ;
      RECT 1165 94415 1415 97945 ;
    LAYER M1 ;
      RECT 1165 98195 1415 99205 ;
    LAYER M1 ;
      RECT 1165 100295 1415 103825 ;
    LAYER M1 ;
      RECT 1165 104075 1415 105085 ;
    LAYER M1 ;
      RECT 1165 106175 1415 109705 ;
    LAYER M1 ;
      RECT 1165 109955 1415 110965 ;
    LAYER M1 ;
      RECT 1165 112055 1415 115585 ;
    LAYER M1 ;
      RECT 1165 115835 1415 116845 ;
    LAYER M1 ;
      RECT 1165 117935 1415 121465 ;
    LAYER M1 ;
      RECT 1165 121715 1415 122725 ;
    LAYER M1 ;
      RECT 1165 123815 1415 127345 ;
    LAYER M1 ;
      RECT 1165 127595 1415 128605 ;
    LAYER M1 ;
      RECT 1165 129695 1415 133225 ;
    LAYER M1 ;
      RECT 1165 133475 1415 134485 ;
    LAYER M1 ;
      RECT 1165 135575 1415 139105 ;
    LAYER M1 ;
      RECT 1165 139355 1415 140365 ;
    LAYER M1 ;
      RECT 1165 141455 1415 144985 ;
    LAYER M1 ;
      RECT 1165 145235 1415 146245 ;
    LAYER M1 ;
      RECT 1165 147335 1415 150865 ;
    LAYER M1 ;
      RECT 1165 151115 1415 152125 ;
    LAYER M1 ;
      RECT 1165 153215 1415 156745 ;
    LAYER M1 ;
      RECT 1165 156995 1415 158005 ;
    LAYER M1 ;
      RECT 1165 159095 1415 162625 ;
    LAYER M1 ;
      RECT 1165 162875 1415 163885 ;
    LAYER M1 ;
      RECT 1165 164975 1415 168505 ;
    LAYER M1 ;
      RECT 1165 168755 1415 169765 ;
    LAYER M1 ;
      RECT 1165 170855 1415 174385 ;
    LAYER M1 ;
      RECT 1165 174635 1415 175645 ;
    LAYER M1 ;
      RECT 1165 176735 1415 180265 ;
    LAYER M1 ;
      RECT 1165 180515 1415 181525 ;
    LAYER M1 ;
      RECT 1165 182615 1415 186145 ;
    LAYER M1 ;
      RECT 1165 186395 1415 187405 ;
    LAYER M1 ;
      RECT 1165 188495 1415 192025 ;
    LAYER M1 ;
      RECT 1165 192275 1415 193285 ;
    LAYER M1 ;
      RECT 1165 194375 1415 197905 ;
    LAYER M1 ;
      RECT 1165 198155 1415 199165 ;
    LAYER M1 ;
      RECT 1165 200255 1415 203785 ;
    LAYER M1 ;
      RECT 1165 204035 1415 205045 ;
    LAYER M1 ;
      RECT 1165 206135 1415 209665 ;
    LAYER M1 ;
      RECT 1165 209915 1415 210925 ;
    LAYER M1 ;
      RECT 1165 212015 1415 215545 ;
    LAYER M1 ;
      RECT 1165 215795 1415 216805 ;
    LAYER M1 ;
      RECT 1165 217895 1415 221425 ;
    LAYER M1 ;
      RECT 1165 221675 1415 222685 ;
    LAYER M1 ;
      RECT 1165 223775 1415 227305 ;
    LAYER M1 ;
      RECT 1165 227555 1415 228565 ;
    LAYER M1 ;
      RECT 1165 229655 1415 233185 ;
    LAYER M1 ;
      RECT 1165 233435 1415 234445 ;
    LAYER M1 ;
      RECT 1165 235535 1415 239065 ;
    LAYER M1 ;
      RECT 1165 239315 1415 240325 ;
    LAYER M1 ;
      RECT 1165 241415 1415 244945 ;
    LAYER M1 ;
      RECT 1165 245195 1415 246205 ;
    LAYER M1 ;
      RECT 1165 247295 1415 250825 ;
    LAYER M1 ;
      RECT 1165 251075 1415 252085 ;
    LAYER M1 ;
      RECT 1165 253175 1415 256705 ;
    LAYER M1 ;
      RECT 1165 256955 1415 257965 ;
    LAYER M1 ;
      RECT 1165 259055 1415 262585 ;
    LAYER M1 ;
      RECT 1165 262835 1415 263845 ;
    LAYER M1 ;
      RECT 1165 264935 1415 268465 ;
    LAYER M1 ;
      RECT 1165 268715 1415 269725 ;
    LAYER M1 ;
      RECT 1165 270815 1415 274345 ;
    LAYER M1 ;
      RECT 1165 274595 1415 275605 ;
    LAYER M1 ;
      RECT 1165 276695 1415 280225 ;
    LAYER M1 ;
      RECT 1165 280475 1415 281485 ;
    LAYER M1 ;
      RECT 1165 282575 1415 286105 ;
    LAYER M1 ;
      RECT 1165 286355 1415 287365 ;
    LAYER M1 ;
      RECT 1165 288455 1415 291985 ;
    LAYER M1 ;
      RECT 1165 292235 1415 293245 ;
    LAYER M1 ;
      RECT 1165 294335 1415 295345 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 735 59135 985 62665 ;
    LAYER M1 ;
      RECT 735 65015 985 68545 ;
    LAYER M1 ;
      RECT 735 70895 985 74425 ;
    LAYER M1 ;
      RECT 735 76775 985 80305 ;
    LAYER M1 ;
      RECT 735 82655 985 86185 ;
    LAYER M1 ;
      RECT 735 88535 985 92065 ;
    LAYER M1 ;
      RECT 735 94415 985 97945 ;
    LAYER M1 ;
      RECT 735 100295 985 103825 ;
    LAYER M1 ;
      RECT 735 106175 985 109705 ;
    LAYER M1 ;
      RECT 735 112055 985 115585 ;
    LAYER M1 ;
      RECT 735 117935 985 121465 ;
    LAYER M1 ;
      RECT 735 123815 985 127345 ;
    LAYER M1 ;
      RECT 735 129695 985 133225 ;
    LAYER M1 ;
      RECT 735 135575 985 139105 ;
    LAYER M1 ;
      RECT 735 141455 985 144985 ;
    LAYER M1 ;
      RECT 735 147335 985 150865 ;
    LAYER M1 ;
      RECT 735 153215 985 156745 ;
    LAYER M1 ;
      RECT 735 159095 985 162625 ;
    LAYER M1 ;
      RECT 735 164975 985 168505 ;
    LAYER M1 ;
      RECT 735 170855 985 174385 ;
    LAYER M1 ;
      RECT 735 176735 985 180265 ;
    LAYER M1 ;
      RECT 735 182615 985 186145 ;
    LAYER M1 ;
      RECT 735 188495 985 192025 ;
    LAYER M1 ;
      RECT 735 194375 985 197905 ;
    LAYER M1 ;
      RECT 735 200255 985 203785 ;
    LAYER M1 ;
      RECT 735 206135 985 209665 ;
    LAYER M1 ;
      RECT 735 212015 985 215545 ;
    LAYER M1 ;
      RECT 735 217895 985 221425 ;
    LAYER M1 ;
      RECT 735 223775 985 227305 ;
    LAYER M1 ;
      RECT 735 229655 985 233185 ;
    LAYER M1 ;
      RECT 735 235535 985 239065 ;
    LAYER M1 ;
      RECT 735 241415 985 244945 ;
    LAYER M1 ;
      RECT 735 247295 985 250825 ;
    LAYER M1 ;
      RECT 735 253175 985 256705 ;
    LAYER M1 ;
      RECT 735 259055 985 262585 ;
    LAYER M1 ;
      RECT 735 264935 985 268465 ;
    LAYER M1 ;
      RECT 735 270815 985 274345 ;
    LAYER M1 ;
      RECT 735 276695 985 280225 ;
    LAYER M1 ;
      RECT 735 282575 985 286105 ;
    LAYER M1 ;
      RECT 735 288455 985 291985 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M1 ;
      RECT 1595 59135 1845 62665 ;
    LAYER M1 ;
      RECT 1595 65015 1845 68545 ;
    LAYER M1 ;
      RECT 1595 70895 1845 74425 ;
    LAYER M1 ;
      RECT 1595 76775 1845 80305 ;
    LAYER M1 ;
      RECT 1595 82655 1845 86185 ;
    LAYER M1 ;
      RECT 1595 88535 1845 92065 ;
    LAYER M1 ;
      RECT 1595 94415 1845 97945 ;
    LAYER M1 ;
      RECT 1595 100295 1845 103825 ;
    LAYER M1 ;
      RECT 1595 106175 1845 109705 ;
    LAYER M1 ;
      RECT 1595 112055 1845 115585 ;
    LAYER M1 ;
      RECT 1595 117935 1845 121465 ;
    LAYER M1 ;
      RECT 1595 123815 1845 127345 ;
    LAYER M1 ;
      RECT 1595 129695 1845 133225 ;
    LAYER M1 ;
      RECT 1595 135575 1845 139105 ;
    LAYER M1 ;
      RECT 1595 141455 1845 144985 ;
    LAYER M1 ;
      RECT 1595 147335 1845 150865 ;
    LAYER M1 ;
      RECT 1595 153215 1845 156745 ;
    LAYER M1 ;
      RECT 1595 159095 1845 162625 ;
    LAYER M1 ;
      RECT 1595 164975 1845 168505 ;
    LAYER M1 ;
      RECT 1595 170855 1845 174385 ;
    LAYER M1 ;
      RECT 1595 176735 1845 180265 ;
    LAYER M1 ;
      RECT 1595 182615 1845 186145 ;
    LAYER M1 ;
      RECT 1595 188495 1845 192025 ;
    LAYER M1 ;
      RECT 1595 194375 1845 197905 ;
    LAYER M1 ;
      RECT 1595 200255 1845 203785 ;
    LAYER M1 ;
      RECT 1595 206135 1845 209665 ;
    LAYER M1 ;
      RECT 1595 212015 1845 215545 ;
    LAYER M1 ;
      RECT 1595 217895 1845 221425 ;
    LAYER M1 ;
      RECT 1595 223775 1845 227305 ;
    LAYER M1 ;
      RECT 1595 229655 1845 233185 ;
    LAYER M1 ;
      RECT 1595 235535 1845 239065 ;
    LAYER M1 ;
      RECT 1595 241415 1845 244945 ;
    LAYER M1 ;
      RECT 1595 247295 1845 250825 ;
    LAYER M1 ;
      RECT 1595 253175 1845 256705 ;
    LAYER M1 ;
      RECT 1595 259055 1845 262585 ;
    LAYER M1 ;
      RECT 1595 264935 1845 268465 ;
    LAYER M1 ;
      RECT 1595 270815 1845 274345 ;
    LAYER M1 ;
      RECT 1595 276695 1845 280225 ;
    LAYER M1 ;
      RECT 1595 282575 1845 286105 ;
    LAYER M1 ;
      RECT 1595 288455 1845 291985 ;
    LAYER M2 ;
      RECT 260 280 1460 560 ;
    LAYER M2 ;
      RECT 260 4480 1460 4760 ;
    LAYER M2 ;
      RECT 690 700 1890 980 ;
    LAYER M2 ;
      RECT 260 6160 1460 6440 ;
    LAYER M2 ;
      RECT 260 10360 1460 10640 ;
    LAYER M2 ;
      RECT 690 6580 1890 6860 ;
    LAYER M2 ;
      RECT 260 12040 1460 12320 ;
    LAYER M2 ;
      RECT 260 16240 1460 16520 ;
    LAYER M2 ;
      RECT 690 12460 1890 12740 ;
    LAYER M2 ;
      RECT 260 17920 1460 18200 ;
    LAYER M2 ;
      RECT 260 22120 1460 22400 ;
    LAYER M2 ;
      RECT 690 18340 1890 18620 ;
    LAYER M2 ;
      RECT 260 23800 1460 24080 ;
    LAYER M2 ;
      RECT 260 28000 1460 28280 ;
    LAYER M2 ;
      RECT 690 24220 1890 24500 ;
    LAYER M2 ;
      RECT 260 29680 1460 29960 ;
    LAYER M2 ;
      RECT 260 33880 1460 34160 ;
    LAYER M2 ;
      RECT 690 30100 1890 30380 ;
    LAYER M2 ;
      RECT 260 35560 1460 35840 ;
    LAYER M2 ;
      RECT 260 39760 1460 40040 ;
    LAYER M2 ;
      RECT 690 35980 1890 36260 ;
    LAYER M2 ;
      RECT 260 41440 1460 41720 ;
    LAYER M2 ;
      RECT 260 45640 1460 45920 ;
    LAYER M2 ;
      RECT 690 41860 1890 42140 ;
    LAYER M2 ;
      RECT 260 47320 1460 47600 ;
    LAYER M2 ;
      RECT 260 51520 1460 51800 ;
    LAYER M2 ;
      RECT 690 47740 1890 48020 ;
    LAYER M2 ;
      RECT 260 53200 1460 53480 ;
    LAYER M2 ;
      RECT 260 57400 1460 57680 ;
    LAYER M2 ;
      RECT 690 53620 1890 53900 ;
    LAYER M2 ;
      RECT 260 59080 1460 59360 ;
    LAYER M2 ;
      RECT 260 63280 1460 63560 ;
    LAYER M2 ;
      RECT 690 59500 1890 59780 ;
    LAYER M2 ;
      RECT 260 64960 1460 65240 ;
    LAYER M2 ;
      RECT 260 69160 1460 69440 ;
    LAYER M2 ;
      RECT 690 65380 1890 65660 ;
    LAYER M2 ;
      RECT 260 70840 1460 71120 ;
    LAYER M2 ;
      RECT 260 75040 1460 75320 ;
    LAYER M2 ;
      RECT 690 71260 1890 71540 ;
    LAYER M2 ;
      RECT 260 76720 1460 77000 ;
    LAYER M2 ;
      RECT 260 80920 1460 81200 ;
    LAYER M2 ;
      RECT 690 77140 1890 77420 ;
    LAYER M2 ;
      RECT 260 82600 1460 82880 ;
    LAYER M2 ;
      RECT 260 86800 1460 87080 ;
    LAYER M2 ;
      RECT 690 83020 1890 83300 ;
    LAYER M2 ;
      RECT 260 88480 1460 88760 ;
    LAYER M2 ;
      RECT 260 92680 1460 92960 ;
    LAYER M2 ;
      RECT 690 88900 1890 89180 ;
    LAYER M2 ;
      RECT 260 94360 1460 94640 ;
    LAYER M2 ;
      RECT 260 98560 1460 98840 ;
    LAYER M2 ;
      RECT 690 94780 1890 95060 ;
    LAYER M2 ;
      RECT 260 100240 1460 100520 ;
    LAYER M2 ;
      RECT 260 104440 1460 104720 ;
    LAYER M2 ;
      RECT 690 100660 1890 100940 ;
    LAYER M2 ;
      RECT 260 106120 1460 106400 ;
    LAYER M2 ;
      RECT 260 110320 1460 110600 ;
    LAYER M2 ;
      RECT 690 106540 1890 106820 ;
    LAYER M2 ;
      RECT 260 112000 1460 112280 ;
    LAYER M2 ;
      RECT 260 116200 1460 116480 ;
    LAYER M2 ;
      RECT 690 112420 1890 112700 ;
    LAYER M2 ;
      RECT 260 117880 1460 118160 ;
    LAYER M2 ;
      RECT 260 122080 1460 122360 ;
    LAYER M2 ;
      RECT 690 118300 1890 118580 ;
    LAYER M2 ;
      RECT 260 123760 1460 124040 ;
    LAYER M2 ;
      RECT 260 127960 1460 128240 ;
    LAYER M2 ;
      RECT 690 124180 1890 124460 ;
    LAYER M2 ;
      RECT 260 129640 1460 129920 ;
    LAYER M2 ;
      RECT 260 133840 1460 134120 ;
    LAYER M2 ;
      RECT 690 130060 1890 130340 ;
    LAYER M2 ;
      RECT 260 135520 1460 135800 ;
    LAYER M2 ;
      RECT 260 139720 1460 140000 ;
    LAYER M2 ;
      RECT 690 135940 1890 136220 ;
    LAYER M2 ;
      RECT 260 141400 1460 141680 ;
    LAYER M2 ;
      RECT 260 145600 1460 145880 ;
    LAYER M2 ;
      RECT 690 141820 1890 142100 ;
    LAYER M2 ;
      RECT 260 147280 1460 147560 ;
    LAYER M2 ;
      RECT 260 151480 1460 151760 ;
    LAYER M2 ;
      RECT 690 147700 1890 147980 ;
    LAYER M2 ;
      RECT 260 153160 1460 153440 ;
    LAYER M2 ;
      RECT 260 157360 1460 157640 ;
    LAYER M2 ;
      RECT 690 153580 1890 153860 ;
    LAYER M2 ;
      RECT 260 159040 1460 159320 ;
    LAYER M2 ;
      RECT 260 163240 1460 163520 ;
    LAYER M2 ;
      RECT 690 159460 1890 159740 ;
    LAYER M2 ;
      RECT 260 164920 1460 165200 ;
    LAYER M2 ;
      RECT 260 169120 1460 169400 ;
    LAYER M2 ;
      RECT 690 165340 1890 165620 ;
    LAYER M2 ;
      RECT 260 170800 1460 171080 ;
    LAYER M2 ;
      RECT 260 175000 1460 175280 ;
    LAYER M2 ;
      RECT 690 171220 1890 171500 ;
    LAYER M2 ;
      RECT 260 176680 1460 176960 ;
    LAYER M2 ;
      RECT 260 180880 1460 181160 ;
    LAYER M2 ;
      RECT 690 177100 1890 177380 ;
    LAYER M2 ;
      RECT 260 182560 1460 182840 ;
    LAYER M2 ;
      RECT 260 186760 1460 187040 ;
    LAYER M2 ;
      RECT 690 182980 1890 183260 ;
    LAYER M2 ;
      RECT 260 188440 1460 188720 ;
    LAYER M2 ;
      RECT 260 192640 1460 192920 ;
    LAYER M2 ;
      RECT 690 188860 1890 189140 ;
    LAYER M2 ;
      RECT 260 194320 1460 194600 ;
    LAYER M2 ;
      RECT 260 198520 1460 198800 ;
    LAYER M2 ;
      RECT 690 194740 1890 195020 ;
    LAYER M2 ;
      RECT 260 200200 1460 200480 ;
    LAYER M2 ;
      RECT 260 204400 1460 204680 ;
    LAYER M2 ;
      RECT 690 200620 1890 200900 ;
    LAYER M2 ;
      RECT 260 206080 1460 206360 ;
    LAYER M2 ;
      RECT 260 210280 1460 210560 ;
    LAYER M2 ;
      RECT 690 206500 1890 206780 ;
    LAYER M2 ;
      RECT 260 211960 1460 212240 ;
    LAYER M2 ;
      RECT 260 216160 1460 216440 ;
    LAYER M2 ;
      RECT 690 212380 1890 212660 ;
    LAYER M2 ;
      RECT 260 217840 1460 218120 ;
    LAYER M2 ;
      RECT 260 222040 1460 222320 ;
    LAYER M2 ;
      RECT 690 218260 1890 218540 ;
    LAYER M2 ;
      RECT 260 223720 1460 224000 ;
    LAYER M2 ;
      RECT 260 227920 1460 228200 ;
    LAYER M2 ;
      RECT 690 224140 1890 224420 ;
    LAYER M2 ;
      RECT 260 229600 1460 229880 ;
    LAYER M2 ;
      RECT 260 233800 1460 234080 ;
    LAYER M2 ;
      RECT 690 230020 1890 230300 ;
    LAYER M2 ;
      RECT 260 235480 1460 235760 ;
    LAYER M2 ;
      RECT 260 239680 1460 239960 ;
    LAYER M2 ;
      RECT 690 235900 1890 236180 ;
    LAYER M2 ;
      RECT 260 241360 1460 241640 ;
    LAYER M2 ;
      RECT 260 245560 1460 245840 ;
    LAYER M2 ;
      RECT 690 241780 1890 242060 ;
    LAYER M2 ;
      RECT 260 247240 1460 247520 ;
    LAYER M2 ;
      RECT 260 251440 1460 251720 ;
    LAYER M2 ;
      RECT 690 247660 1890 247940 ;
    LAYER M2 ;
      RECT 260 253120 1460 253400 ;
    LAYER M2 ;
      RECT 260 257320 1460 257600 ;
    LAYER M2 ;
      RECT 690 253540 1890 253820 ;
    LAYER M2 ;
      RECT 260 259000 1460 259280 ;
    LAYER M2 ;
      RECT 260 263200 1460 263480 ;
    LAYER M2 ;
      RECT 690 259420 1890 259700 ;
    LAYER M2 ;
      RECT 260 264880 1460 265160 ;
    LAYER M2 ;
      RECT 260 269080 1460 269360 ;
    LAYER M2 ;
      RECT 690 265300 1890 265580 ;
    LAYER M2 ;
      RECT 260 270760 1460 271040 ;
    LAYER M2 ;
      RECT 260 274960 1460 275240 ;
    LAYER M2 ;
      RECT 690 271180 1890 271460 ;
    LAYER M2 ;
      RECT 260 276640 1460 276920 ;
    LAYER M2 ;
      RECT 260 280840 1460 281120 ;
    LAYER M2 ;
      RECT 690 277060 1890 277340 ;
    LAYER M2 ;
      RECT 260 282520 1460 282800 ;
    LAYER M2 ;
      RECT 260 286720 1460 287000 ;
    LAYER M2 ;
      RECT 690 282940 1890 283220 ;
    LAYER M2 ;
      RECT 260 288400 1460 288680 ;
    LAYER M2 ;
      RECT 260 292600 1460 292880 ;
    LAYER M2 ;
      RECT 690 294700 1890 294980 ;
    LAYER M2 ;
      RECT 690 288820 1890 289100 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53255 1375 53425 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59135 1375 59305 ;
    LAYER V1 ;
      RECT 1205 63335 1375 63505 ;
    LAYER V1 ;
      RECT 1205 65015 1375 65185 ;
    LAYER V1 ;
      RECT 1205 69215 1375 69385 ;
    LAYER V1 ;
      RECT 1205 70895 1375 71065 ;
    LAYER V1 ;
      RECT 1205 75095 1375 75265 ;
    LAYER V1 ;
      RECT 1205 76775 1375 76945 ;
    LAYER V1 ;
      RECT 1205 80975 1375 81145 ;
    LAYER V1 ;
      RECT 1205 82655 1375 82825 ;
    LAYER V1 ;
      RECT 1205 86855 1375 87025 ;
    LAYER V1 ;
      RECT 1205 88535 1375 88705 ;
    LAYER V1 ;
      RECT 1205 92735 1375 92905 ;
    LAYER V1 ;
      RECT 1205 94415 1375 94585 ;
    LAYER V1 ;
      RECT 1205 98615 1375 98785 ;
    LAYER V1 ;
      RECT 1205 100295 1375 100465 ;
    LAYER V1 ;
      RECT 1205 104495 1375 104665 ;
    LAYER V1 ;
      RECT 1205 106175 1375 106345 ;
    LAYER V1 ;
      RECT 1205 110375 1375 110545 ;
    LAYER V1 ;
      RECT 1205 112055 1375 112225 ;
    LAYER V1 ;
      RECT 1205 116255 1375 116425 ;
    LAYER V1 ;
      RECT 1205 117935 1375 118105 ;
    LAYER V1 ;
      RECT 1205 122135 1375 122305 ;
    LAYER V1 ;
      RECT 1205 123815 1375 123985 ;
    LAYER V1 ;
      RECT 1205 128015 1375 128185 ;
    LAYER V1 ;
      RECT 1205 129695 1375 129865 ;
    LAYER V1 ;
      RECT 1205 133895 1375 134065 ;
    LAYER V1 ;
      RECT 1205 135575 1375 135745 ;
    LAYER V1 ;
      RECT 1205 139775 1375 139945 ;
    LAYER V1 ;
      RECT 1205 141455 1375 141625 ;
    LAYER V1 ;
      RECT 1205 145655 1375 145825 ;
    LAYER V1 ;
      RECT 1205 147335 1375 147505 ;
    LAYER V1 ;
      RECT 1205 151535 1375 151705 ;
    LAYER V1 ;
      RECT 1205 153215 1375 153385 ;
    LAYER V1 ;
      RECT 1205 157415 1375 157585 ;
    LAYER V1 ;
      RECT 1205 159095 1375 159265 ;
    LAYER V1 ;
      RECT 1205 163295 1375 163465 ;
    LAYER V1 ;
      RECT 1205 164975 1375 165145 ;
    LAYER V1 ;
      RECT 1205 169175 1375 169345 ;
    LAYER V1 ;
      RECT 1205 170855 1375 171025 ;
    LAYER V1 ;
      RECT 1205 175055 1375 175225 ;
    LAYER V1 ;
      RECT 1205 176735 1375 176905 ;
    LAYER V1 ;
      RECT 1205 180935 1375 181105 ;
    LAYER V1 ;
      RECT 1205 182615 1375 182785 ;
    LAYER V1 ;
      RECT 1205 186815 1375 186985 ;
    LAYER V1 ;
      RECT 1205 188495 1375 188665 ;
    LAYER V1 ;
      RECT 1205 192695 1375 192865 ;
    LAYER V1 ;
      RECT 1205 194375 1375 194545 ;
    LAYER V1 ;
      RECT 1205 198575 1375 198745 ;
    LAYER V1 ;
      RECT 1205 200255 1375 200425 ;
    LAYER V1 ;
      RECT 1205 204455 1375 204625 ;
    LAYER V1 ;
      RECT 1205 206135 1375 206305 ;
    LAYER V1 ;
      RECT 1205 210335 1375 210505 ;
    LAYER V1 ;
      RECT 1205 212015 1375 212185 ;
    LAYER V1 ;
      RECT 1205 216215 1375 216385 ;
    LAYER V1 ;
      RECT 1205 217895 1375 218065 ;
    LAYER V1 ;
      RECT 1205 222095 1375 222265 ;
    LAYER V1 ;
      RECT 1205 223775 1375 223945 ;
    LAYER V1 ;
      RECT 1205 227975 1375 228145 ;
    LAYER V1 ;
      RECT 1205 229655 1375 229825 ;
    LAYER V1 ;
      RECT 1205 233855 1375 234025 ;
    LAYER V1 ;
      RECT 1205 235535 1375 235705 ;
    LAYER V1 ;
      RECT 1205 239735 1375 239905 ;
    LAYER V1 ;
      RECT 1205 241415 1375 241585 ;
    LAYER V1 ;
      RECT 1205 245615 1375 245785 ;
    LAYER V1 ;
      RECT 1205 247295 1375 247465 ;
    LAYER V1 ;
      RECT 1205 251495 1375 251665 ;
    LAYER V1 ;
      RECT 1205 253175 1375 253345 ;
    LAYER V1 ;
      RECT 1205 257375 1375 257545 ;
    LAYER V1 ;
      RECT 1205 259055 1375 259225 ;
    LAYER V1 ;
      RECT 1205 263255 1375 263425 ;
    LAYER V1 ;
      RECT 1205 264935 1375 265105 ;
    LAYER V1 ;
      RECT 1205 269135 1375 269305 ;
    LAYER V1 ;
      RECT 1205 270815 1375 270985 ;
    LAYER V1 ;
      RECT 1205 275015 1375 275185 ;
    LAYER V1 ;
      RECT 1205 276695 1375 276865 ;
    LAYER V1 ;
      RECT 1205 280895 1375 281065 ;
    LAYER V1 ;
      RECT 1205 282575 1375 282745 ;
    LAYER V1 ;
      RECT 1205 286775 1375 286945 ;
    LAYER V1 ;
      RECT 1205 288455 1375 288625 ;
    LAYER V1 ;
      RECT 1205 292655 1375 292825 ;
    LAYER V1 ;
      RECT 1205 294755 1375 294925 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 775 53675 945 53845 ;
    LAYER V1 ;
      RECT 775 59555 945 59725 ;
    LAYER V1 ;
      RECT 775 65435 945 65605 ;
    LAYER V1 ;
      RECT 775 71315 945 71485 ;
    LAYER V1 ;
      RECT 775 77195 945 77365 ;
    LAYER V1 ;
      RECT 775 83075 945 83245 ;
    LAYER V1 ;
      RECT 775 88955 945 89125 ;
    LAYER V1 ;
      RECT 775 94835 945 95005 ;
    LAYER V1 ;
      RECT 775 100715 945 100885 ;
    LAYER V1 ;
      RECT 775 106595 945 106765 ;
    LAYER V1 ;
      RECT 775 112475 945 112645 ;
    LAYER V1 ;
      RECT 775 118355 945 118525 ;
    LAYER V1 ;
      RECT 775 124235 945 124405 ;
    LAYER V1 ;
      RECT 775 130115 945 130285 ;
    LAYER V1 ;
      RECT 775 135995 945 136165 ;
    LAYER V1 ;
      RECT 775 141875 945 142045 ;
    LAYER V1 ;
      RECT 775 147755 945 147925 ;
    LAYER V1 ;
      RECT 775 153635 945 153805 ;
    LAYER V1 ;
      RECT 775 159515 945 159685 ;
    LAYER V1 ;
      RECT 775 165395 945 165565 ;
    LAYER V1 ;
      RECT 775 171275 945 171445 ;
    LAYER V1 ;
      RECT 775 177155 945 177325 ;
    LAYER V1 ;
      RECT 775 183035 945 183205 ;
    LAYER V1 ;
      RECT 775 188915 945 189085 ;
    LAYER V1 ;
      RECT 775 194795 945 194965 ;
    LAYER V1 ;
      RECT 775 200675 945 200845 ;
    LAYER V1 ;
      RECT 775 206555 945 206725 ;
    LAYER V1 ;
      RECT 775 212435 945 212605 ;
    LAYER V1 ;
      RECT 775 218315 945 218485 ;
    LAYER V1 ;
      RECT 775 224195 945 224365 ;
    LAYER V1 ;
      RECT 775 230075 945 230245 ;
    LAYER V1 ;
      RECT 775 235955 945 236125 ;
    LAYER V1 ;
      RECT 775 241835 945 242005 ;
    LAYER V1 ;
      RECT 775 247715 945 247885 ;
    LAYER V1 ;
      RECT 775 253595 945 253765 ;
    LAYER V1 ;
      RECT 775 259475 945 259645 ;
    LAYER V1 ;
      RECT 775 265355 945 265525 ;
    LAYER V1 ;
      RECT 775 271235 945 271405 ;
    LAYER V1 ;
      RECT 775 277115 945 277285 ;
    LAYER V1 ;
      RECT 775 282995 945 283165 ;
    LAYER V1 ;
      RECT 775 288875 945 289045 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 1635 53675 1805 53845 ;
    LAYER V1 ;
      RECT 1635 59555 1805 59725 ;
    LAYER V1 ;
      RECT 1635 65435 1805 65605 ;
    LAYER V1 ;
      RECT 1635 71315 1805 71485 ;
    LAYER V1 ;
      RECT 1635 77195 1805 77365 ;
    LAYER V1 ;
      RECT 1635 83075 1805 83245 ;
    LAYER V1 ;
      RECT 1635 88955 1805 89125 ;
    LAYER V1 ;
      RECT 1635 94835 1805 95005 ;
    LAYER V1 ;
      RECT 1635 100715 1805 100885 ;
    LAYER V1 ;
      RECT 1635 106595 1805 106765 ;
    LAYER V1 ;
      RECT 1635 112475 1805 112645 ;
    LAYER V1 ;
      RECT 1635 118355 1805 118525 ;
    LAYER V1 ;
      RECT 1635 124235 1805 124405 ;
    LAYER V1 ;
      RECT 1635 130115 1805 130285 ;
    LAYER V1 ;
      RECT 1635 135995 1805 136165 ;
    LAYER V1 ;
      RECT 1635 141875 1805 142045 ;
    LAYER V1 ;
      RECT 1635 147755 1805 147925 ;
    LAYER V1 ;
      RECT 1635 153635 1805 153805 ;
    LAYER V1 ;
      RECT 1635 159515 1805 159685 ;
    LAYER V1 ;
      RECT 1635 165395 1805 165565 ;
    LAYER V1 ;
      RECT 1635 171275 1805 171445 ;
    LAYER V1 ;
      RECT 1635 177155 1805 177325 ;
    LAYER V1 ;
      RECT 1635 183035 1805 183205 ;
    LAYER V1 ;
      RECT 1635 188915 1805 189085 ;
    LAYER V1 ;
      RECT 1635 194795 1805 194965 ;
    LAYER V1 ;
      RECT 1635 200675 1805 200845 ;
    LAYER V1 ;
      RECT 1635 206555 1805 206725 ;
    LAYER V1 ;
      RECT 1635 212435 1805 212605 ;
    LAYER V1 ;
      RECT 1635 218315 1805 218485 ;
    LAYER V1 ;
      RECT 1635 224195 1805 224365 ;
    LAYER V1 ;
      RECT 1635 230075 1805 230245 ;
    LAYER V1 ;
      RECT 1635 235955 1805 236125 ;
    LAYER V1 ;
      RECT 1635 241835 1805 242005 ;
    LAYER V1 ;
      RECT 1635 247715 1805 247885 ;
    LAYER V1 ;
      RECT 1635 253595 1805 253765 ;
    LAYER V1 ;
      RECT 1635 259475 1805 259645 ;
    LAYER V1 ;
      RECT 1635 265355 1805 265525 ;
    LAYER V1 ;
      RECT 1635 271235 1805 271405 ;
    LAYER V1 ;
      RECT 1635 277115 1805 277285 ;
    LAYER V1 ;
      RECT 1635 282995 1805 283165 ;
    LAYER V1 ;
      RECT 1635 288875 1805 289045 ;
    LAYER V2 ;
      RECT 1215 345 1365 495 ;
    LAYER V2 ;
      RECT 1215 4545 1365 4695 ;
    LAYER V2 ;
      RECT 1215 6225 1365 6375 ;
    LAYER V2 ;
      RECT 1215 10425 1365 10575 ;
    LAYER V2 ;
      RECT 1215 12105 1365 12255 ;
    LAYER V2 ;
      RECT 1215 16305 1365 16455 ;
    LAYER V2 ;
      RECT 1215 17985 1365 18135 ;
    LAYER V2 ;
      RECT 1215 22185 1365 22335 ;
    LAYER V2 ;
      RECT 1215 23865 1365 24015 ;
    LAYER V2 ;
      RECT 1215 28065 1365 28215 ;
    LAYER V2 ;
      RECT 1215 29745 1365 29895 ;
    LAYER V2 ;
      RECT 1215 33945 1365 34095 ;
    LAYER V2 ;
      RECT 1215 35625 1365 35775 ;
    LAYER V2 ;
      RECT 1215 39825 1365 39975 ;
    LAYER V2 ;
      RECT 1215 41505 1365 41655 ;
    LAYER V2 ;
      RECT 1215 45705 1365 45855 ;
    LAYER V2 ;
      RECT 1215 47385 1365 47535 ;
    LAYER V2 ;
      RECT 1215 51585 1365 51735 ;
    LAYER V2 ;
      RECT 1215 53265 1365 53415 ;
    LAYER V2 ;
      RECT 1215 57465 1365 57615 ;
    LAYER V2 ;
      RECT 1215 59145 1365 59295 ;
    LAYER V2 ;
      RECT 1215 63345 1365 63495 ;
    LAYER V2 ;
      RECT 1215 65025 1365 65175 ;
    LAYER V2 ;
      RECT 1215 69225 1365 69375 ;
    LAYER V2 ;
      RECT 1215 70905 1365 71055 ;
    LAYER V2 ;
      RECT 1215 75105 1365 75255 ;
    LAYER V2 ;
      RECT 1215 76785 1365 76935 ;
    LAYER V2 ;
      RECT 1215 80985 1365 81135 ;
    LAYER V2 ;
      RECT 1215 82665 1365 82815 ;
    LAYER V2 ;
      RECT 1215 86865 1365 87015 ;
    LAYER V2 ;
      RECT 1215 88545 1365 88695 ;
    LAYER V2 ;
      RECT 1215 92745 1365 92895 ;
    LAYER V2 ;
      RECT 1215 94425 1365 94575 ;
    LAYER V2 ;
      RECT 1215 98625 1365 98775 ;
    LAYER V2 ;
      RECT 1215 100305 1365 100455 ;
    LAYER V2 ;
      RECT 1215 104505 1365 104655 ;
    LAYER V2 ;
      RECT 1215 106185 1365 106335 ;
    LAYER V2 ;
      RECT 1215 110385 1365 110535 ;
    LAYER V2 ;
      RECT 1215 112065 1365 112215 ;
    LAYER V2 ;
      RECT 1215 116265 1365 116415 ;
    LAYER V2 ;
      RECT 1215 117945 1365 118095 ;
    LAYER V2 ;
      RECT 1215 122145 1365 122295 ;
    LAYER V2 ;
      RECT 1215 123825 1365 123975 ;
    LAYER V2 ;
      RECT 1215 128025 1365 128175 ;
    LAYER V2 ;
      RECT 1215 129705 1365 129855 ;
    LAYER V2 ;
      RECT 1215 133905 1365 134055 ;
    LAYER V2 ;
      RECT 1215 135585 1365 135735 ;
    LAYER V2 ;
      RECT 1215 139785 1365 139935 ;
    LAYER V2 ;
      RECT 1215 141465 1365 141615 ;
    LAYER V2 ;
      RECT 1215 145665 1365 145815 ;
    LAYER V2 ;
      RECT 1215 147345 1365 147495 ;
    LAYER V2 ;
      RECT 1215 151545 1365 151695 ;
    LAYER V2 ;
      RECT 1215 153225 1365 153375 ;
    LAYER V2 ;
      RECT 1215 157425 1365 157575 ;
    LAYER V2 ;
      RECT 1215 159105 1365 159255 ;
    LAYER V2 ;
      RECT 1215 163305 1365 163455 ;
    LAYER V2 ;
      RECT 1215 164985 1365 165135 ;
    LAYER V2 ;
      RECT 1215 169185 1365 169335 ;
    LAYER V2 ;
      RECT 1215 170865 1365 171015 ;
    LAYER V2 ;
      RECT 1215 175065 1365 175215 ;
    LAYER V2 ;
      RECT 1215 176745 1365 176895 ;
    LAYER V2 ;
      RECT 1215 180945 1365 181095 ;
    LAYER V2 ;
      RECT 1215 182625 1365 182775 ;
    LAYER V2 ;
      RECT 1215 186825 1365 186975 ;
    LAYER V2 ;
      RECT 1215 188505 1365 188655 ;
    LAYER V2 ;
      RECT 1215 192705 1365 192855 ;
    LAYER V2 ;
      RECT 1215 194385 1365 194535 ;
    LAYER V2 ;
      RECT 1215 198585 1365 198735 ;
    LAYER V2 ;
      RECT 1215 200265 1365 200415 ;
    LAYER V2 ;
      RECT 1215 204465 1365 204615 ;
    LAYER V2 ;
      RECT 1215 206145 1365 206295 ;
    LAYER V2 ;
      RECT 1215 210345 1365 210495 ;
    LAYER V2 ;
      RECT 1215 212025 1365 212175 ;
    LAYER V2 ;
      RECT 1215 216225 1365 216375 ;
    LAYER V2 ;
      RECT 1215 217905 1365 218055 ;
    LAYER V2 ;
      RECT 1215 222105 1365 222255 ;
    LAYER V2 ;
      RECT 1215 223785 1365 223935 ;
    LAYER V2 ;
      RECT 1215 227985 1365 228135 ;
    LAYER V2 ;
      RECT 1215 229665 1365 229815 ;
    LAYER V2 ;
      RECT 1215 233865 1365 234015 ;
    LAYER V2 ;
      RECT 1215 235545 1365 235695 ;
    LAYER V2 ;
      RECT 1215 239745 1365 239895 ;
    LAYER V2 ;
      RECT 1215 241425 1365 241575 ;
    LAYER V2 ;
      RECT 1215 245625 1365 245775 ;
    LAYER V2 ;
      RECT 1215 247305 1365 247455 ;
    LAYER V2 ;
      RECT 1215 251505 1365 251655 ;
    LAYER V2 ;
      RECT 1215 253185 1365 253335 ;
    LAYER V2 ;
      RECT 1215 257385 1365 257535 ;
    LAYER V2 ;
      RECT 1215 259065 1365 259215 ;
    LAYER V2 ;
      RECT 1215 263265 1365 263415 ;
    LAYER V2 ;
      RECT 1215 264945 1365 265095 ;
    LAYER V2 ;
      RECT 1215 269145 1365 269295 ;
    LAYER V2 ;
      RECT 1215 270825 1365 270975 ;
    LAYER V2 ;
      RECT 1215 275025 1365 275175 ;
    LAYER V2 ;
      RECT 1215 276705 1365 276855 ;
    LAYER V2 ;
      RECT 1215 280905 1365 281055 ;
    LAYER V2 ;
      RECT 1215 282585 1365 282735 ;
    LAYER V2 ;
      RECT 1215 286785 1365 286935 ;
    LAYER V2 ;
      RECT 1215 288465 1365 288615 ;
    LAYER V2 ;
      RECT 1215 292665 1365 292815 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 6645 1795 6795 ;
    LAYER V2 ;
      RECT 1645 12525 1795 12675 ;
    LAYER V2 ;
      RECT 1645 18405 1795 18555 ;
    LAYER V2 ;
      RECT 1645 24285 1795 24435 ;
    LAYER V2 ;
      RECT 1645 30165 1795 30315 ;
    LAYER V2 ;
      RECT 1645 36045 1795 36195 ;
    LAYER V2 ;
      RECT 1645 41925 1795 42075 ;
    LAYER V2 ;
      RECT 1645 47805 1795 47955 ;
    LAYER V2 ;
      RECT 1645 53685 1795 53835 ;
    LAYER V2 ;
      RECT 1645 59565 1795 59715 ;
    LAYER V2 ;
      RECT 1645 65445 1795 65595 ;
    LAYER V2 ;
      RECT 1645 71325 1795 71475 ;
    LAYER V2 ;
      RECT 1645 77205 1795 77355 ;
    LAYER V2 ;
      RECT 1645 83085 1795 83235 ;
    LAYER V2 ;
      RECT 1645 88965 1795 89115 ;
    LAYER V2 ;
      RECT 1645 94845 1795 94995 ;
    LAYER V2 ;
      RECT 1645 100725 1795 100875 ;
    LAYER V2 ;
      RECT 1645 106605 1795 106755 ;
    LAYER V2 ;
      RECT 1645 112485 1795 112635 ;
    LAYER V2 ;
      RECT 1645 118365 1795 118515 ;
    LAYER V2 ;
      RECT 1645 124245 1795 124395 ;
    LAYER V2 ;
      RECT 1645 130125 1795 130275 ;
    LAYER V2 ;
      RECT 1645 136005 1795 136155 ;
    LAYER V2 ;
      RECT 1645 141885 1795 142035 ;
    LAYER V2 ;
      RECT 1645 147765 1795 147915 ;
    LAYER V2 ;
      RECT 1645 153645 1795 153795 ;
    LAYER V2 ;
      RECT 1645 159525 1795 159675 ;
    LAYER V2 ;
      RECT 1645 165405 1795 165555 ;
    LAYER V2 ;
      RECT 1645 171285 1795 171435 ;
    LAYER V2 ;
      RECT 1645 177165 1795 177315 ;
    LAYER V2 ;
      RECT 1645 183045 1795 183195 ;
    LAYER V2 ;
      RECT 1645 188925 1795 189075 ;
    LAYER V2 ;
      RECT 1645 194805 1795 194955 ;
    LAYER V2 ;
      RECT 1645 200685 1795 200835 ;
    LAYER V2 ;
      RECT 1645 206565 1795 206715 ;
    LAYER V2 ;
      RECT 1645 212445 1795 212595 ;
    LAYER V2 ;
      RECT 1645 218325 1795 218475 ;
    LAYER V2 ;
      RECT 1645 224205 1795 224355 ;
    LAYER V2 ;
      RECT 1645 230085 1795 230235 ;
    LAYER V2 ;
      RECT 1645 235965 1795 236115 ;
    LAYER V2 ;
      RECT 1645 241845 1795 241995 ;
    LAYER V2 ;
      RECT 1645 247725 1795 247875 ;
    LAYER V2 ;
      RECT 1645 253605 1795 253755 ;
    LAYER V2 ;
      RECT 1645 259485 1795 259635 ;
    LAYER V2 ;
      RECT 1645 265365 1795 265515 ;
    LAYER V2 ;
      RECT 1645 271245 1795 271395 ;
    LAYER V2 ;
      RECT 1645 277125 1795 277275 ;
    LAYER V2 ;
      RECT 1645 283005 1795 283155 ;
    LAYER V2 ;
      RECT 1645 288885 1795 289035 ;
    LAYER V2 ;
      RECT 1645 294765 1795 294915 ;
  END
END DCL_NMOS_S_38019457_X1_Y50
